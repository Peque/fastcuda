


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Librabry for instantiating Xilinx primitives
Library UNISIM;
use UNISIM.vcomponents.all;

-- Library for using arithmetic functions with signed/unsigned values
use IEEE.NUMERIC_STD.ALL;




entity smem is
end smem;

architecture Behavioral of smem is

begin

BRAM_TDP_MACRO_inst : BRAM_TDP_MACRO

generic map (

	-- Memory size and target device family
	BRAM_SIZE => "9Kb",
	DEVICE => "SPARTAN6",

	-- Optional port output register
	DOA_REG => 0,
	DOB_REG => 0,

	-- Initial values on ports
	INIT_A => X"000000000",
	INIT_B => X"000000000",
	INIT_FILE => "NONE",

	-- Read and write width (must be equal)
	READ_WIDTH_A  => 32,
	WRITE_WIDTH_A => 32,
	READ_WIDTH_B  => 32,
	WRITE_WIDTH_B => 32,

	-- Warning produced and affected outputs/memory location go unknown
	SIM_COLLISION_CHECK => "ALL",

	-- Output value on the DO ports upon the assertion of the syncronous reset signal
	SRVAL_A => X"000000000",
	SRVAL_B => X"000000000",

	-- NO_CHANGE mode: the output latches remain unchanged during a write operation
	WRITE_MODE_A => "NO_CHANGE",
	WRITE_MODE_B => "NO_CHANGE",

	-- Initial contents of the RAM
	INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

	-- Parity bits initialization
	INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"

) port map (

	DOA => DOA,        -- Output port-A data
	DOB => DOB,        -- Output port-B data
	ADDRA => ADDRA,    -- Input port-A address
	ADDRB => ADDRB,    -- Input port-B address
	CLKA => CLKA,      -- Input port-A clock
	CLKB => CLKB,      -- Input port-B clock
	DIA => DIA,        -- Input port-A data
	DIB => DIB,        -- Input port-B data
	ENA => ENA,        -- Input port-A enable
	ENB => ENB,        -- Input port-B enable
	REGCEA => REGCEA,  -- Input port-A output register enable
	REGCEB => REGCEB,  -- Input port-B output register enable
	RSTA => RSTA,      -- Input port-A reset
	RSTB => RSTB,      -- Input port-B reset
	WEA => WEA,        -- Input port-A write enable
	WEB => WEB         -- Input port-B write enable

);

end Behavioral;

