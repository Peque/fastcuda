--
-- smem.vhd
--
-- Copyright 2012 Miguel Sánchez de León Peque <msdeleonpeque@gmail.com>
--
-- This program is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program; if not, write to the Free Software
-- Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston,
-- MA 02110-1301, USA.
--
--



library ieee;
use ieee.std_logic_1164.all;

library unisim;
use unisim.vcomponents.all;

library unimacro;
use unimacro.vcomponents.all;



entity smem is

	generic (

		N_PORTS         : integer := 32;
		N_BRAMS         : integer := 16;
		LOG2_N_PORTS    : integer := 5  -- TODO: should be calculated from N_PORTS and then used only to generate the VHDL code

	);

	port (

		DO                     : out std_logic_vector(32 * N_PORTS - 1 downto 0);    -- Data output ports
		DI                     : in  std_logic_vector(32 * N_PORTS - 1 downto 0);    -- Data input ports
		ADDR_0, ADDR_1, ADDR_2, ADDR_3, ADDR_4, ADDR_5, ADDR_6, ADDR_7, ADDR_8, ADDR_9, ADDR_10, ADDR_11, ADDR_12, ADDR_13, ADDR_14, ADDR_15, ADDR_16, ADDR_17, ADDR_18, ADDR_19, ADDR_20, ADDR_21, ADDR_22, ADDR_23, ADDR_24, ADDR_25, ADDR_26, ADDR_27, ADDR_28, ADDR_29, ADDR_30, ADDR_31     : in  std_logic_vector(12 downto 0);    -- Address input ports
		WE_0, WE_1, WE_2, WE_3, WE_4, WE_5, WE_6, WE_7, WE_8, WE_9, WE_10, WE_11, WE_12, WE_13, WE_14, WE_15, WE_16, WE_17, WE_18, WE_19, WE_20, WE_21, WE_22, WE_23, WE_24, WE_25, WE_26, WE_27, WE_28, WE_29, WE_30, WE_31                     : in  std_logic_vector(3 downto 0);     -- Byte write enable input ports
		BRAM_CLK, TRIG_CLK, RST                                            : in  std_logic;                        -- Clock and reset input ports
		REQ_0, REQ_1, REQ_2, REQ_3, REQ_4, REQ_5, REQ_6, REQ_7, REQ_8, REQ_9, REQ_10, REQ_11, REQ_12, REQ_13, REQ_14, REQ_15, REQ_16, REQ_17, REQ_18, REQ_19, REQ_20, REQ_21, REQ_22, REQ_23, REQ_24, REQ_25, REQ_26, REQ_27, REQ_28, REQ_29, REQ_30, REQ_31             : in  std_logic;                        -- Request input ports
		RDY_0, RDY_1, RDY_2, RDY_3, RDY_4, RDY_5, RDY_6, RDY_7, RDY_8, RDY_9, RDY_10, RDY_11, RDY_12, RDY_13, RDY_14, RDY_15, RDY_16, RDY_17, RDY_18, RDY_19, RDY_20, RDY_21, RDY_22, RDY_23, RDY_24, RDY_25, RDY_26, RDY_27, RDY_28, RDY_29, RDY_30, RDY_31             : out std_logic                         -- Ready output port

	);

end smem;



architecture smem_arch of smem is


	constant DIP_value         : std_logic_vector(3 downto 0) := "0000";
	constant LOWADDR_value     : std_logic_vector(4 downto 0) := "00000";
	constant REGCE_value       : std_logic := '0';
	constant EN_value          : std_logic := '1';

	signal k0_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k1_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k2_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k3_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k4_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k5_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k6_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k7_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k8_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k9_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k10_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k11_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k12_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k13_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k14_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k15_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k16_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k17_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k18_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k19_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k20_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k21_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k22_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k23_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k24_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k25_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k26_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k27_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k28_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k29_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k30_output_sel       : bit_vector(4 downto 0) := "00000";
	signal k31_output_sel       : bit_vector(4 downto 0) := "00000";

	signal k0_being_served     : bit := '0';
	signal k1_being_served     : bit := '0';
	signal k2_being_served     : bit := '0';
	signal k3_being_served     : bit := '0';
	signal k4_being_served     : bit := '0';
	signal k5_being_served     : bit := '0';
	signal k6_being_served     : bit := '0';
	signal k7_being_served     : bit := '0';
	signal k8_being_served     : bit := '0';
	signal k9_being_served     : bit := '0';
	signal k10_being_served     : bit := '0';
	signal k11_being_served     : bit := '0';
	signal k12_being_served     : bit := '0';
	signal k13_being_served     : bit := '0';
	signal k14_being_served     : bit := '0';
	signal k15_being_served     : bit := '0';
	signal k16_being_served     : bit := '0';
	signal k17_being_served     : bit := '0';
	signal k18_being_served     : bit := '0';
	signal k19_being_served     : bit := '0';
	signal k20_being_served     : bit := '0';
	signal k21_being_served     : bit := '0';
	signal k22_being_served     : bit := '0';
	signal k23_being_served     : bit := '0';
	signal k24_being_served     : bit := '0';
	signal k25_being_served     : bit := '0';
	signal k26_being_served     : bit := '0';
	signal k27_being_served     : bit := '0';
	signal k28_being_served     : bit := '0';
	signal k29_being_served     : bit := '0';
	signal k30_being_served     : bit := '0';
	signal k31_being_served     : bit := '0';

	signal k0_needs_attention  : bit := '0';
	signal k1_needs_attention  : bit := '0';
	signal k2_needs_attention  : bit := '0';
	signal k3_needs_attention  : bit := '0';
	signal k4_needs_attention  : bit := '0';
	signal k5_needs_attention  : bit := '0';
	signal k6_needs_attention  : bit := '0';
	signal k7_needs_attention  : bit := '0';
	signal k8_needs_attention  : bit := '0';
	signal k9_needs_attention  : bit := '0';
	signal k10_needs_attention  : bit := '0';
	signal k11_needs_attention  : bit := '0';
	signal k12_needs_attention  : bit := '0';
	signal k13_needs_attention  : bit := '0';
	signal k14_needs_attention  : bit := '0';
	signal k15_needs_attention  : bit := '0';
	signal k16_needs_attention  : bit := '0';
	signal k17_needs_attention  : bit := '0';
	signal k18_needs_attention  : bit := '0';
	signal k19_needs_attention  : bit := '0';
	signal k20_needs_attention  : bit := '0';
	signal k21_needs_attention  : bit := '0';
	signal k22_needs_attention  : bit := '0';
	signal k23_needs_attention  : bit := '0';
	signal k24_needs_attention  : bit := '0';
	signal k25_needs_attention  : bit := '0';
	signal k26_needs_attention  : bit := '0';
	signal k27_needs_attention  : bit := '0';
	signal k28_needs_attention  : bit := '0';
	signal k29_needs_attention  : bit := '0';
	signal k30_needs_attention  : bit := '0';
	signal k31_needs_attention  : bit := '0';

	signal addr_0_eq_addr_1    : bit := '0';
	signal addr_0_eq_addr_2    : bit := '0';
	signal addr_0_eq_addr_3    : bit := '0';
	signal addr_0_eq_addr_4    : bit := '0';
	signal addr_0_eq_addr_5    : bit := '0';
	signal addr_0_eq_addr_6    : bit := '0';
	signal addr_0_eq_addr_7    : bit := '0';
	signal addr_0_eq_addr_8    : bit := '0';
	signal addr_0_eq_addr_9    : bit := '0';
	signal addr_0_eq_addr_10    : bit := '0';
	signal addr_0_eq_addr_11    : bit := '0';
	signal addr_0_eq_addr_12    : bit := '0';
	signal addr_0_eq_addr_13    : bit := '0';
	signal addr_0_eq_addr_14    : bit := '0';
	signal addr_0_eq_addr_15    : bit := '0';
	signal addr_0_eq_addr_16    : bit := '0';
	signal addr_0_eq_addr_17    : bit := '0';
	signal addr_0_eq_addr_18    : bit := '0';
	signal addr_0_eq_addr_19    : bit := '0';
	signal addr_0_eq_addr_20    : bit := '0';
	signal addr_0_eq_addr_21    : bit := '0';
	signal addr_0_eq_addr_22    : bit := '0';
	signal addr_0_eq_addr_23    : bit := '0';
	signal addr_0_eq_addr_24    : bit := '0';
	signal addr_0_eq_addr_25    : bit := '0';
	signal addr_0_eq_addr_26    : bit := '0';
	signal addr_0_eq_addr_27    : bit := '0';
	signal addr_0_eq_addr_28    : bit := '0';
	signal addr_0_eq_addr_29    : bit := '0';
	signal addr_0_eq_addr_30    : bit := '0';
	signal addr_0_eq_addr_31    : bit := '0';
	signal addr_1_eq_addr_2    : bit := '0';
	signal addr_1_eq_addr_3    : bit := '0';
	signal addr_1_eq_addr_4    : bit := '0';
	signal addr_1_eq_addr_5    : bit := '0';
	signal addr_1_eq_addr_6    : bit := '0';
	signal addr_1_eq_addr_7    : bit := '0';
	signal addr_1_eq_addr_8    : bit := '0';
	signal addr_1_eq_addr_9    : bit := '0';
	signal addr_1_eq_addr_10    : bit := '0';
	signal addr_1_eq_addr_11    : bit := '0';
	signal addr_1_eq_addr_12    : bit := '0';
	signal addr_1_eq_addr_13    : bit := '0';
	signal addr_1_eq_addr_14    : bit := '0';
	signal addr_1_eq_addr_15    : bit := '0';
	signal addr_1_eq_addr_16    : bit := '0';
	signal addr_1_eq_addr_17    : bit := '0';
	signal addr_1_eq_addr_18    : bit := '0';
	signal addr_1_eq_addr_19    : bit := '0';
	signal addr_1_eq_addr_20    : bit := '0';
	signal addr_1_eq_addr_21    : bit := '0';
	signal addr_1_eq_addr_22    : bit := '0';
	signal addr_1_eq_addr_23    : bit := '0';
	signal addr_1_eq_addr_24    : bit := '0';
	signal addr_1_eq_addr_25    : bit := '0';
	signal addr_1_eq_addr_26    : bit := '0';
	signal addr_1_eq_addr_27    : bit := '0';
	signal addr_1_eq_addr_28    : bit := '0';
	signal addr_1_eq_addr_29    : bit := '0';
	signal addr_1_eq_addr_30    : bit := '0';
	signal addr_1_eq_addr_31    : bit := '0';
	signal addr_2_eq_addr_3    : bit := '0';
	signal addr_2_eq_addr_4    : bit := '0';
	signal addr_2_eq_addr_5    : bit := '0';
	signal addr_2_eq_addr_6    : bit := '0';
	signal addr_2_eq_addr_7    : bit := '0';
	signal addr_2_eq_addr_8    : bit := '0';
	signal addr_2_eq_addr_9    : bit := '0';
	signal addr_2_eq_addr_10    : bit := '0';
	signal addr_2_eq_addr_11    : bit := '0';
	signal addr_2_eq_addr_12    : bit := '0';
	signal addr_2_eq_addr_13    : bit := '0';
	signal addr_2_eq_addr_14    : bit := '0';
	signal addr_2_eq_addr_15    : bit := '0';
	signal addr_2_eq_addr_16    : bit := '0';
	signal addr_2_eq_addr_17    : bit := '0';
	signal addr_2_eq_addr_18    : bit := '0';
	signal addr_2_eq_addr_19    : bit := '0';
	signal addr_2_eq_addr_20    : bit := '0';
	signal addr_2_eq_addr_21    : bit := '0';
	signal addr_2_eq_addr_22    : bit := '0';
	signal addr_2_eq_addr_23    : bit := '0';
	signal addr_2_eq_addr_24    : bit := '0';
	signal addr_2_eq_addr_25    : bit := '0';
	signal addr_2_eq_addr_26    : bit := '0';
	signal addr_2_eq_addr_27    : bit := '0';
	signal addr_2_eq_addr_28    : bit := '0';
	signal addr_2_eq_addr_29    : bit := '0';
	signal addr_2_eq_addr_30    : bit := '0';
	signal addr_2_eq_addr_31    : bit := '0';
	signal addr_3_eq_addr_4    : bit := '0';
	signal addr_3_eq_addr_5    : bit := '0';
	signal addr_3_eq_addr_6    : bit := '0';
	signal addr_3_eq_addr_7    : bit := '0';
	signal addr_3_eq_addr_8    : bit := '0';
	signal addr_3_eq_addr_9    : bit := '0';
	signal addr_3_eq_addr_10    : bit := '0';
	signal addr_3_eq_addr_11    : bit := '0';
	signal addr_3_eq_addr_12    : bit := '0';
	signal addr_3_eq_addr_13    : bit := '0';
	signal addr_3_eq_addr_14    : bit := '0';
	signal addr_3_eq_addr_15    : bit := '0';
	signal addr_3_eq_addr_16    : bit := '0';
	signal addr_3_eq_addr_17    : bit := '0';
	signal addr_3_eq_addr_18    : bit := '0';
	signal addr_3_eq_addr_19    : bit := '0';
	signal addr_3_eq_addr_20    : bit := '0';
	signal addr_3_eq_addr_21    : bit := '0';
	signal addr_3_eq_addr_22    : bit := '0';
	signal addr_3_eq_addr_23    : bit := '0';
	signal addr_3_eq_addr_24    : bit := '0';
	signal addr_3_eq_addr_25    : bit := '0';
	signal addr_3_eq_addr_26    : bit := '0';
	signal addr_3_eq_addr_27    : bit := '0';
	signal addr_3_eq_addr_28    : bit := '0';
	signal addr_3_eq_addr_29    : bit := '0';
	signal addr_3_eq_addr_30    : bit := '0';
	signal addr_3_eq_addr_31    : bit := '0';
	signal addr_4_eq_addr_5    : bit := '0';
	signal addr_4_eq_addr_6    : bit := '0';
	signal addr_4_eq_addr_7    : bit := '0';
	signal addr_4_eq_addr_8    : bit := '0';
	signal addr_4_eq_addr_9    : bit := '0';
	signal addr_4_eq_addr_10    : bit := '0';
	signal addr_4_eq_addr_11    : bit := '0';
	signal addr_4_eq_addr_12    : bit := '0';
	signal addr_4_eq_addr_13    : bit := '0';
	signal addr_4_eq_addr_14    : bit := '0';
	signal addr_4_eq_addr_15    : bit := '0';
	signal addr_4_eq_addr_16    : bit := '0';
	signal addr_4_eq_addr_17    : bit := '0';
	signal addr_4_eq_addr_18    : bit := '0';
	signal addr_4_eq_addr_19    : bit := '0';
	signal addr_4_eq_addr_20    : bit := '0';
	signal addr_4_eq_addr_21    : bit := '0';
	signal addr_4_eq_addr_22    : bit := '0';
	signal addr_4_eq_addr_23    : bit := '0';
	signal addr_4_eq_addr_24    : bit := '0';
	signal addr_4_eq_addr_25    : bit := '0';
	signal addr_4_eq_addr_26    : bit := '0';
	signal addr_4_eq_addr_27    : bit := '0';
	signal addr_4_eq_addr_28    : bit := '0';
	signal addr_4_eq_addr_29    : bit := '0';
	signal addr_4_eq_addr_30    : bit := '0';
	signal addr_4_eq_addr_31    : bit := '0';
	signal addr_5_eq_addr_6    : bit := '0';
	signal addr_5_eq_addr_7    : bit := '0';
	signal addr_5_eq_addr_8    : bit := '0';
	signal addr_5_eq_addr_9    : bit := '0';
	signal addr_5_eq_addr_10    : bit := '0';
	signal addr_5_eq_addr_11    : bit := '0';
	signal addr_5_eq_addr_12    : bit := '0';
	signal addr_5_eq_addr_13    : bit := '0';
	signal addr_5_eq_addr_14    : bit := '0';
	signal addr_5_eq_addr_15    : bit := '0';
	signal addr_5_eq_addr_16    : bit := '0';
	signal addr_5_eq_addr_17    : bit := '0';
	signal addr_5_eq_addr_18    : bit := '0';
	signal addr_5_eq_addr_19    : bit := '0';
	signal addr_5_eq_addr_20    : bit := '0';
	signal addr_5_eq_addr_21    : bit := '0';
	signal addr_5_eq_addr_22    : bit := '0';
	signal addr_5_eq_addr_23    : bit := '0';
	signal addr_5_eq_addr_24    : bit := '0';
	signal addr_5_eq_addr_25    : bit := '0';
	signal addr_5_eq_addr_26    : bit := '0';
	signal addr_5_eq_addr_27    : bit := '0';
	signal addr_5_eq_addr_28    : bit := '0';
	signal addr_5_eq_addr_29    : bit := '0';
	signal addr_5_eq_addr_30    : bit := '0';
	signal addr_5_eq_addr_31    : bit := '0';
	signal addr_6_eq_addr_7    : bit := '0';
	signal addr_6_eq_addr_8    : bit := '0';
	signal addr_6_eq_addr_9    : bit := '0';
	signal addr_6_eq_addr_10    : bit := '0';
	signal addr_6_eq_addr_11    : bit := '0';
	signal addr_6_eq_addr_12    : bit := '0';
	signal addr_6_eq_addr_13    : bit := '0';
	signal addr_6_eq_addr_14    : bit := '0';
	signal addr_6_eq_addr_15    : bit := '0';
	signal addr_6_eq_addr_16    : bit := '0';
	signal addr_6_eq_addr_17    : bit := '0';
	signal addr_6_eq_addr_18    : bit := '0';
	signal addr_6_eq_addr_19    : bit := '0';
	signal addr_6_eq_addr_20    : bit := '0';
	signal addr_6_eq_addr_21    : bit := '0';
	signal addr_6_eq_addr_22    : bit := '0';
	signal addr_6_eq_addr_23    : bit := '0';
	signal addr_6_eq_addr_24    : bit := '0';
	signal addr_6_eq_addr_25    : bit := '0';
	signal addr_6_eq_addr_26    : bit := '0';
	signal addr_6_eq_addr_27    : bit := '0';
	signal addr_6_eq_addr_28    : bit := '0';
	signal addr_6_eq_addr_29    : bit := '0';
	signal addr_6_eq_addr_30    : bit := '0';
	signal addr_6_eq_addr_31    : bit := '0';
	signal addr_7_eq_addr_8    : bit := '0';
	signal addr_7_eq_addr_9    : bit := '0';
	signal addr_7_eq_addr_10    : bit := '0';
	signal addr_7_eq_addr_11    : bit := '0';
	signal addr_7_eq_addr_12    : bit := '0';
	signal addr_7_eq_addr_13    : bit := '0';
	signal addr_7_eq_addr_14    : bit := '0';
	signal addr_7_eq_addr_15    : bit := '0';
	signal addr_7_eq_addr_16    : bit := '0';
	signal addr_7_eq_addr_17    : bit := '0';
	signal addr_7_eq_addr_18    : bit := '0';
	signal addr_7_eq_addr_19    : bit := '0';
	signal addr_7_eq_addr_20    : bit := '0';
	signal addr_7_eq_addr_21    : bit := '0';
	signal addr_7_eq_addr_22    : bit := '0';
	signal addr_7_eq_addr_23    : bit := '0';
	signal addr_7_eq_addr_24    : bit := '0';
	signal addr_7_eq_addr_25    : bit := '0';
	signal addr_7_eq_addr_26    : bit := '0';
	signal addr_7_eq_addr_27    : bit := '0';
	signal addr_7_eq_addr_28    : bit := '0';
	signal addr_7_eq_addr_29    : bit := '0';
	signal addr_7_eq_addr_30    : bit := '0';
	signal addr_7_eq_addr_31    : bit := '0';
	signal addr_8_eq_addr_9    : bit := '0';
	signal addr_8_eq_addr_10    : bit := '0';
	signal addr_8_eq_addr_11    : bit := '0';
	signal addr_8_eq_addr_12    : bit := '0';
	signal addr_8_eq_addr_13    : bit := '0';
	signal addr_8_eq_addr_14    : bit := '0';
	signal addr_8_eq_addr_15    : bit := '0';
	signal addr_8_eq_addr_16    : bit := '0';
	signal addr_8_eq_addr_17    : bit := '0';
	signal addr_8_eq_addr_18    : bit := '0';
	signal addr_8_eq_addr_19    : bit := '0';
	signal addr_8_eq_addr_20    : bit := '0';
	signal addr_8_eq_addr_21    : bit := '0';
	signal addr_8_eq_addr_22    : bit := '0';
	signal addr_8_eq_addr_23    : bit := '0';
	signal addr_8_eq_addr_24    : bit := '0';
	signal addr_8_eq_addr_25    : bit := '0';
	signal addr_8_eq_addr_26    : bit := '0';
	signal addr_8_eq_addr_27    : bit := '0';
	signal addr_8_eq_addr_28    : bit := '0';
	signal addr_8_eq_addr_29    : bit := '0';
	signal addr_8_eq_addr_30    : bit := '0';
	signal addr_8_eq_addr_31    : bit := '0';
	signal addr_9_eq_addr_10    : bit := '0';
	signal addr_9_eq_addr_11    : bit := '0';
	signal addr_9_eq_addr_12    : bit := '0';
	signal addr_9_eq_addr_13    : bit := '0';
	signal addr_9_eq_addr_14    : bit := '0';
	signal addr_9_eq_addr_15    : bit := '0';
	signal addr_9_eq_addr_16    : bit := '0';
	signal addr_9_eq_addr_17    : bit := '0';
	signal addr_9_eq_addr_18    : bit := '0';
	signal addr_9_eq_addr_19    : bit := '0';
	signal addr_9_eq_addr_20    : bit := '0';
	signal addr_9_eq_addr_21    : bit := '0';
	signal addr_9_eq_addr_22    : bit := '0';
	signal addr_9_eq_addr_23    : bit := '0';
	signal addr_9_eq_addr_24    : bit := '0';
	signal addr_9_eq_addr_25    : bit := '0';
	signal addr_9_eq_addr_26    : bit := '0';
	signal addr_9_eq_addr_27    : bit := '0';
	signal addr_9_eq_addr_28    : bit := '0';
	signal addr_9_eq_addr_29    : bit := '0';
	signal addr_9_eq_addr_30    : bit := '0';
	signal addr_9_eq_addr_31    : bit := '0';
	signal addr_10_eq_addr_11    : bit := '0';
	signal addr_10_eq_addr_12    : bit := '0';
	signal addr_10_eq_addr_13    : bit := '0';
	signal addr_10_eq_addr_14    : bit := '0';
	signal addr_10_eq_addr_15    : bit := '0';
	signal addr_10_eq_addr_16    : bit := '0';
	signal addr_10_eq_addr_17    : bit := '0';
	signal addr_10_eq_addr_18    : bit := '0';
	signal addr_10_eq_addr_19    : bit := '0';
	signal addr_10_eq_addr_20    : bit := '0';
	signal addr_10_eq_addr_21    : bit := '0';
	signal addr_10_eq_addr_22    : bit := '0';
	signal addr_10_eq_addr_23    : bit := '0';
	signal addr_10_eq_addr_24    : bit := '0';
	signal addr_10_eq_addr_25    : bit := '0';
	signal addr_10_eq_addr_26    : bit := '0';
	signal addr_10_eq_addr_27    : bit := '0';
	signal addr_10_eq_addr_28    : bit := '0';
	signal addr_10_eq_addr_29    : bit := '0';
	signal addr_10_eq_addr_30    : bit := '0';
	signal addr_10_eq_addr_31    : bit := '0';
	signal addr_11_eq_addr_12    : bit := '0';
	signal addr_11_eq_addr_13    : bit := '0';
	signal addr_11_eq_addr_14    : bit := '0';
	signal addr_11_eq_addr_15    : bit := '0';
	signal addr_11_eq_addr_16    : bit := '0';
	signal addr_11_eq_addr_17    : bit := '0';
	signal addr_11_eq_addr_18    : bit := '0';
	signal addr_11_eq_addr_19    : bit := '0';
	signal addr_11_eq_addr_20    : bit := '0';
	signal addr_11_eq_addr_21    : bit := '0';
	signal addr_11_eq_addr_22    : bit := '0';
	signal addr_11_eq_addr_23    : bit := '0';
	signal addr_11_eq_addr_24    : bit := '0';
	signal addr_11_eq_addr_25    : bit := '0';
	signal addr_11_eq_addr_26    : bit := '0';
	signal addr_11_eq_addr_27    : bit := '0';
	signal addr_11_eq_addr_28    : bit := '0';
	signal addr_11_eq_addr_29    : bit := '0';
	signal addr_11_eq_addr_30    : bit := '0';
	signal addr_11_eq_addr_31    : bit := '0';
	signal addr_12_eq_addr_13    : bit := '0';
	signal addr_12_eq_addr_14    : bit := '0';
	signal addr_12_eq_addr_15    : bit := '0';
	signal addr_12_eq_addr_16    : bit := '0';
	signal addr_12_eq_addr_17    : bit := '0';
	signal addr_12_eq_addr_18    : bit := '0';
	signal addr_12_eq_addr_19    : bit := '0';
	signal addr_12_eq_addr_20    : bit := '0';
	signal addr_12_eq_addr_21    : bit := '0';
	signal addr_12_eq_addr_22    : bit := '0';
	signal addr_12_eq_addr_23    : bit := '0';
	signal addr_12_eq_addr_24    : bit := '0';
	signal addr_12_eq_addr_25    : bit := '0';
	signal addr_12_eq_addr_26    : bit := '0';
	signal addr_12_eq_addr_27    : bit := '0';
	signal addr_12_eq_addr_28    : bit := '0';
	signal addr_12_eq_addr_29    : bit := '0';
	signal addr_12_eq_addr_30    : bit := '0';
	signal addr_12_eq_addr_31    : bit := '0';
	signal addr_13_eq_addr_14    : bit := '0';
	signal addr_13_eq_addr_15    : bit := '0';
	signal addr_13_eq_addr_16    : bit := '0';
	signal addr_13_eq_addr_17    : bit := '0';
	signal addr_13_eq_addr_18    : bit := '0';
	signal addr_13_eq_addr_19    : bit := '0';
	signal addr_13_eq_addr_20    : bit := '0';
	signal addr_13_eq_addr_21    : bit := '0';
	signal addr_13_eq_addr_22    : bit := '0';
	signal addr_13_eq_addr_23    : bit := '0';
	signal addr_13_eq_addr_24    : bit := '0';
	signal addr_13_eq_addr_25    : bit := '0';
	signal addr_13_eq_addr_26    : bit := '0';
	signal addr_13_eq_addr_27    : bit := '0';
	signal addr_13_eq_addr_28    : bit := '0';
	signal addr_13_eq_addr_29    : bit := '0';
	signal addr_13_eq_addr_30    : bit := '0';
	signal addr_13_eq_addr_31    : bit := '0';
	signal addr_14_eq_addr_15    : bit := '0';
	signal addr_14_eq_addr_16    : bit := '0';
	signal addr_14_eq_addr_17    : bit := '0';
	signal addr_14_eq_addr_18    : bit := '0';
	signal addr_14_eq_addr_19    : bit := '0';
	signal addr_14_eq_addr_20    : bit := '0';
	signal addr_14_eq_addr_21    : bit := '0';
	signal addr_14_eq_addr_22    : bit := '0';
	signal addr_14_eq_addr_23    : bit := '0';
	signal addr_14_eq_addr_24    : bit := '0';
	signal addr_14_eq_addr_25    : bit := '0';
	signal addr_14_eq_addr_26    : bit := '0';
	signal addr_14_eq_addr_27    : bit := '0';
	signal addr_14_eq_addr_28    : bit := '0';
	signal addr_14_eq_addr_29    : bit := '0';
	signal addr_14_eq_addr_30    : bit := '0';
	signal addr_14_eq_addr_31    : bit := '0';
	signal addr_15_eq_addr_16    : bit := '0';
	signal addr_15_eq_addr_17    : bit := '0';
	signal addr_15_eq_addr_18    : bit := '0';
	signal addr_15_eq_addr_19    : bit := '0';
	signal addr_15_eq_addr_20    : bit := '0';
	signal addr_15_eq_addr_21    : bit := '0';
	signal addr_15_eq_addr_22    : bit := '0';
	signal addr_15_eq_addr_23    : bit := '0';
	signal addr_15_eq_addr_24    : bit := '0';
	signal addr_15_eq_addr_25    : bit := '0';
	signal addr_15_eq_addr_26    : bit := '0';
	signal addr_15_eq_addr_27    : bit := '0';
	signal addr_15_eq_addr_28    : bit := '0';
	signal addr_15_eq_addr_29    : bit := '0';
	signal addr_15_eq_addr_30    : bit := '0';
	signal addr_15_eq_addr_31    : bit := '0';
	signal addr_16_eq_addr_17    : bit := '0';
	signal addr_16_eq_addr_18    : bit := '0';
	signal addr_16_eq_addr_19    : bit := '0';
	signal addr_16_eq_addr_20    : bit := '0';
	signal addr_16_eq_addr_21    : bit := '0';
	signal addr_16_eq_addr_22    : bit := '0';
	signal addr_16_eq_addr_23    : bit := '0';
	signal addr_16_eq_addr_24    : bit := '0';
	signal addr_16_eq_addr_25    : bit := '0';
	signal addr_16_eq_addr_26    : bit := '0';
	signal addr_16_eq_addr_27    : bit := '0';
	signal addr_16_eq_addr_28    : bit := '0';
	signal addr_16_eq_addr_29    : bit := '0';
	signal addr_16_eq_addr_30    : bit := '0';
	signal addr_16_eq_addr_31    : bit := '0';
	signal addr_17_eq_addr_18    : bit := '0';
	signal addr_17_eq_addr_19    : bit := '0';
	signal addr_17_eq_addr_20    : bit := '0';
	signal addr_17_eq_addr_21    : bit := '0';
	signal addr_17_eq_addr_22    : bit := '0';
	signal addr_17_eq_addr_23    : bit := '0';
	signal addr_17_eq_addr_24    : bit := '0';
	signal addr_17_eq_addr_25    : bit := '0';
	signal addr_17_eq_addr_26    : bit := '0';
	signal addr_17_eq_addr_27    : bit := '0';
	signal addr_17_eq_addr_28    : bit := '0';
	signal addr_17_eq_addr_29    : bit := '0';
	signal addr_17_eq_addr_30    : bit := '0';
	signal addr_17_eq_addr_31    : bit := '0';
	signal addr_18_eq_addr_19    : bit := '0';
	signal addr_18_eq_addr_20    : bit := '0';
	signal addr_18_eq_addr_21    : bit := '0';
	signal addr_18_eq_addr_22    : bit := '0';
	signal addr_18_eq_addr_23    : bit := '0';
	signal addr_18_eq_addr_24    : bit := '0';
	signal addr_18_eq_addr_25    : bit := '0';
	signal addr_18_eq_addr_26    : bit := '0';
	signal addr_18_eq_addr_27    : bit := '0';
	signal addr_18_eq_addr_28    : bit := '0';
	signal addr_18_eq_addr_29    : bit := '0';
	signal addr_18_eq_addr_30    : bit := '0';
	signal addr_18_eq_addr_31    : bit := '0';
	signal addr_19_eq_addr_20    : bit := '0';
	signal addr_19_eq_addr_21    : bit := '0';
	signal addr_19_eq_addr_22    : bit := '0';
	signal addr_19_eq_addr_23    : bit := '0';
	signal addr_19_eq_addr_24    : bit := '0';
	signal addr_19_eq_addr_25    : bit := '0';
	signal addr_19_eq_addr_26    : bit := '0';
	signal addr_19_eq_addr_27    : bit := '0';
	signal addr_19_eq_addr_28    : bit := '0';
	signal addr_19_eq_addr_29    : bit := '0';
	signal addr_19_eq_addr_30    : bit := '0';
	signal addr_19_eq_addr_31    : bit := '0';
	signal addr_20_eq_addr_21    : bit := '0';
	signal addr_20_eq_addr_22    : bit := '0';
	signal addr_20_eq_addr_23    : bit := '0';
	signal addr_20_eq_addr_24    : bit := '0';
	signal addr_20_eq_addr_25    : bit := '0';
	signal addr_20_eq_addr_26    : bit := '0';
	signal addr_20_eq_addr_27    : bit := '0';
	signal addr_20_eq_addr_28    : bit := '0';
	signal addr_20_eq_addr_29    : bit := '0';
	signal addr_20_eq_addr_30    : bit := '0';
	signal addr_20_eq_addr_31    : bit := '0';
	signal addr_21_eq_addr_22    : bit := '0';
	signal addr_21_eq_addr_23    : bit := '0';
	signal addr_21_eq_addr_24    : bit := '0';
	signal addr_21_eq_addr_25    : bit := '0';
	signal addr_21_eq_addr_26    : bit := '0';
	signal addr_21_eq_addr_27    : bit := '0';
	signal addr_21_eq_addr_28    : bit := '0';
	signal addr_21_eq_addr_29    : bit := '0';
	signal addr_21_eq_addr_30    : bit := '0';
	signal addr_21_eq_addr_31    : bit := '0';
	signal addr_22_eq_addr_23    : bit := '0';
	signal addr_22_eq_addr_24    : bit := '0';
	signal addr_22_eq_addr_25    : bit := '0';
	signal addr_22_eq_addr_26    : bit := '0';
	signal addr_22_eq_addr_27    : bit := '0';
	signal addr_22_eq_addr_28    : bit := '0';
	signal addr_22_eq_addr_29    : bit := '0';
	signal addr_22_eq_addr_30    : bit := '0';
	signal addr_22_eq_addr_31    : bit := '0';
	signal addr_23_eq_addr_24    : bit := '0';
	signal addr_23_eq_addr_25    : bit := '0';
	signal addr_23_eq_addr_26    : bit := '0';
	signal addr_23_eq_addr_27    : bit := '0';
	signal addr_23_eq_addr_28    : bit := '0';
	signal addr_23_eq_addr_29    : bit := '0';
	signal addr_23_eq_addr_30    : bit := '0';
	signal addr_23_eq_addr_31    : bit := '0';
	signal addr_24_eq_addr_25    : bit := '0';
	signal addr_24_eq_addr_26    : bit := '0';
	signal addr_24_eq_addr_27    : bit := '0';
	signal addr_24_eq_addr_28    : bit := '0';
	signal addr_24_eq_addr_29    : bit := '0';
	signal addr_24_eq_addr_30    : bit := '0';
	signal addr_24_eq_addr_31    : bit := '0';
	signal addr_25_eq_addr_26    : bit := '0';
	signal addr_25_eq_addr_27    : bit := '0';
	signal addr_25_eq_addr_28    : bit := '0';
	signal addr_25_eq_addr_29    : bit := '0';
	signal addr_25_eq_addr_30    : bit := '0';
	signal addr_25_eq_addr_31    : bit := '0';
	signal addr_26_eq_addr_27    : bit := '0';
	signal addr_26_eq_addr_28    : bit := '0';
	signal addr_26_eq_addr_29    : bit := '0';
	signal addr_26_eq_addr_30    : bit := '0';
	signal addr_26_eq_addr_31    : bit := '0';
	signal addr_27_eq_addr_28    : bit := '0';
	signal addr_27_eq_addr_29    : bit := '0';
	signal addr_27_eq_addr_30    : bit := '0';
	signal addr_27_eq_addr_31    : bit := '0';
	signal addr_28_eq_addr_29    : bit := '0';
	signal addr_28_eq_addr_30    : bit := '0';
	signal addr_28_eq_addr_31    : bit := '0';
	signal addr_29_eq_addr_30    : bit := '0';
	signal addr_29_eq_addr_31    : bit := '0';
	signal addr_30_eq_addr_31    : bit := '0';

	signal we_0_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_1_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_2_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_3_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_4_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_5_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_6_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_7_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_8_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_9_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_10_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_11_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_12_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_13_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_14_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_15_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_16_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_17_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_18_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_19_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_20_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_21_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_22_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_23_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_24_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_25_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_26_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_27_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_28_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_29_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_30_safe           : std_logic_vector(3 downto 0) := "0000";
	signal we_31_safe           : std_logic_vector(3 downto 0) := "0000";

	signal bram_0_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_1_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_2_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_3_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_4_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_5_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_6_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_7_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_8_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_9_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_10_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_11_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_12_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_13_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_14_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_15_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_16_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_17_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_18_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_19_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_20_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_21_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_22_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_23_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_24_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_25_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_26_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_27_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_28_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_29_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_30_input_sel    : bit_vector(4 downto 0) := "00000";
	signal bram_31_input_sel    : bit_vector(4 downto 0) := "00000";

	signal k0_needs_bram_0     : bit := '0';
	signal k0_needs_bram_1     : bit := '0';
	signal k0_needs_bram_2     : bit := '0';
	signal k0_needs_bram_3     : bit := '0';
	signal k0_needs_bram_4     : bit := '0';
	signal k0_needs_bram_5     : bit := '0';
	signal k0_needs_bram_6     : bit := '0';
	signal k0_needs_bram_7     : bit := '0';
	signal k0_needs_bram_8     : bit := '0';
	signal k0_needs_bram_9     : bit := '0';
	signal k0_needs_bram_10     : bit := '0';
	signal k0_needs_bram_11     : bit := '0';
	signal k0_needs_bram_12     : bit := '0';
	signal k0_needs_bram_13     : bit := '0';
	signal k0_needs_bram_14     : bit := '0';
	signal k0_needs_bram_15     : bit := '0';
	signal k1_needs_bram_0     : bit := '0';
	signal k1_needs_bram_1     : bit := '0';
	signal k1_needs_bram_2     : bit := '0';
	signal k1_needs_bram_3     : bit := '0';
	signal k1_needs_bram_4     : bit := '0';
	signal k1_needs_bram_5     : bit := '0';
	signal k1_needs_bram_6     : bit := '0';
	signal k1_needs_bram_7     : bit := '0';
	signal k1_needs_bram_8     : bit := '0';
	signal k1_needs_bram_9     : bit := '0';
	signal k1_needs_bram_10     : bit := '0';
	signal k1_needs_bram_11     : bit := '0';
	signal k1_needs_bram_12     : bit := '0';
	signal k1_needs_bram_13     : bit := '0';
	signal k1_needs_bram_14     : bit := '0';
	signal k1_needs_bram_15     : bit := '0';
	signal k2_needs_bram_0     : bit := '0';
	signal k2_needs_bram_1     : bit := '0';
	signal k2_needs_bram_2     : bit := '0';
	signal k2_needs_bram_3     : bit := '0';
	signal k2_needs_bram_4     : bit := '0';
	signal k2_needs_bram_5     : bit := '0';
	signal k2_needs_bram_6     : bit := '0';
	signal k2_needs_bram_7     : bit := '0';
	signal k2_needs_bram_8     : bit := '0';
	signal k2_needs_bram_9     : bit := '0';
	signal k2_needs_bram_10     : bit := '0';
	signal k2_needs_bram_11     : bit := '0';
	signal k2_needs_bram_12     : bit := '0';
	signal k2_needs_bram_13     : bit := '0';
	signal k2_needs_bram_14     : bit := '0';
	signal k2_needs_bram_15     : bit := '0';
	signal k3_needs_bram_0     : bit := '0';
	signal k3_needs_bram_1     : bit := '0';
	signal k3_needs_bram_2     : bit := '0';
	signal k3_needs_bram_3     : bit := '0';
	signal k3_needs_bram_4     : bit := '0';
	signal k3_needs_bram_5     : bit := '0';
	signal k3_needs_bram_6     : bit := '0';
	signal k3_needs_bram_7     : bit := '0';
	signal k3_needs_bram_8     : bit := '0';
	signal k3_needs_bram_9     : bit := '0';
	signal k3_needs_bram_10     : bit := '0';
	signal k3_needs_bram_11     : bit := '0';
	signal k3_needs_bram_12     : bit := '0';
	signal k3_needs_bram_13     : bit := '0';
	signal k3_needs_bram_14     : bit := '0';
	signal k3_needs_bram_15     : bit := '0';
	signal k4_needs_bram_0     : bit := '0';
	signal k4_needs_bram_1     : bit := '0';
	signal k4_needs_bram_2     : bit := '0';
	signal k4_needs_bram_3     : bit := '0';
	signal k4_needs_bram_4     : bit := '0';
	signal k4_needs_bram_5     : bit := '0';
	signal k4_needs_bram_6     : bit := '0';
	signal k4_needs_bram_7     : bit := '0';
	signal k4_needs_bram_8     : bit := '0';
	signal k4_needs_bram_9     : bit := '0';
	signal k4_needs_bram_10     : bit := '0';
	signal k4_needs_bram_11     : bit := '0';
	signal k4_needs_bram_12     : bit := '0';
	signal k4_needs_bram_13     : bit := '0';
	signal k4_needs_bram_14     : bit := '0';
	signal k4_needs_bram_15     : bit := '0';
	signal k5_needs_bram_0     : bit := '0';
	signal k5_needs_bram_1     : bit := '0';
	signal k5_needs_bram_2     : bit := '0';
	signal k5_needs_bram_3     : bit := '0';
	signal k5_needs_bram_4     : bit := '0';
	signal k5_needs_bram_5     : bit := '0';
	signal k5_needs_bram_6     : bit := '0';
	signal k5_needs_bram_7     : bit := '0';
	signal k5_needs_bram_8     : bit := '0';
	signal k5_needs_bram_9     : bit := '0';
	signal k5_needs_bram_10     : bit := '0';
	signal k5_needs_bram_11     : bit := '0';
	signal k5_needs_bram_12     : bit := '0';
	signal k5_needs_bram_13     : bit := '0';
	signal k5_needs_bram_14     : bit := '0';
	signal k5_needs_bram_15     : bit := '0';
	signal k6_needs_bram_0     : bit := '0';
	signal k6_needs_bram_1     : bit := '0';
	signal k6_needs_bram_2     : bit := '0';
	signal k6_needs_bram_3     : bit := '0';
	signal k6_needs_bram_4     : bit := '0';
	signal k6_needs_bram_5     : bit := '0';
	signal k6_needs_bram_6     : bit := '0';
	signal k6_needs_bram_7     : bit := '0';
	signal k6_needs_bram_8     : bit := '0';
	signal k6_needs_bram_9     : bit := '0';
	signal k6_needs_bram_10     : bit := '0';
	signal k6_needs_bram_11     : bit := '0';
	signal k6_needs_bram_12     : bit := '0';
	signal k6_needs_bram_13     : bit := '0';
	signal k6_needs_bram_14     : bit := '0';
	signal k6_needs_bram_15     : bit := '0';
	signal k7_needs_bram_0     : bit := '0';
	signal k7_needs_bram_1     : bit := '0';
	signal k7_needs_bram_2     : bit := '0';
	signal k7_needs_bram_3     : bit := '0';
	signal k7_needs_bram_4     : bit := '0';
	signal k7_needs_bram_5     : bit := '0';
	signal k7_needs_bram_6     : bit := '0';
	signal k7_needs_bram_7     : bit := '0';
	signal k7_needs_bram_8     : bit := '0';
	signal k7_needs_bram_9     : bit := '0';
	signal k7_needs_bram_10     : bit := '0';
	signal k7_needs_bram_11     : bit := '0';
	signal k7_needs_bram_12     : bit := '0';
	signal k7_needs_bram_13     : bit := '0';
	signal k7_needs_bram_14     : bit := '0';
	signal k7_needs_bram_15     : bit := '0';
	signal k8_needs_bram_0     : bit := '0';
	signal k8_needs_bram_1     : bit := '0';
	signal k8_needs_bram_2     : bit := '0';
	signal k8_needs_bram_3     : bit := '0';
	signal k8_needs_bram_4     : bit := '0';
	signal k8_needs_bram_5     : bit := '0';
	signal k8_needs_bram_6     : bit := '0';
	signal k8_needs_bram_7     : bit := '0';
	signal k8_needs_bram_8     : bit := '0';
	signal k8_needs_bram_9     : bit := '0';
	signal k8_needs_bram_10     : bit := '0';
	signal k8_needs_bram_11     : bit := '0';
	signal k8_needs_bram_12     : bit := '0';
	signal k8_needs_bram_13     : bit := '0';
	signal k8_needs_bram_14     : bit := '0';
	signal k8_needs_bram_15     : bit := '0';
	signal k9_needs_bram_0     : bit := '0';
	signal k9_needs_bram_1     : bit := '0';
	signal k9_needs_bram_2     : bit := '0';
	signal k9_needs_bram_3     : bit := '0';
	signal k9_needs_bram_4     : bit := '0';
	signal k9_needs_bram_5     : bit := '0';
	signal k9_needs_bram_6     : bit := '0';
	signal k9_needs_bram_7     : bit := '0';
	signal k9_needs_bram_8     : bit := '0';
	signal k9_needs_bram_9     : bit := '0';
	signal k9_needs_bram_10     : bit := '0';
	signal k9_needs_bram_11     : bit := '0';
	signal k9_needs_bram_12     : bit := '0';
	signal k9_needs_bram_13     : bit := '0';
	signal k9_needs_bram_14     : bit := '0';
	signal k9_needs_bram_15     : bit := '0';
	signal k10_needs_bram_0     : bit := '0';
	signal k10_needs_bram_1     : bit := '0';
	signal k10_needs_bram_2     : bit := '0';
	signal k10_needs_bram_3     : bit := '0';
	signal k10_needs_bram_4     : bit := '0';
	signal k10_needs_bram_5     : bit := '0';
	signal k10_needs_bram_6     : bit := '0';
	signal k10_needs_bram_7     : bit := '0';
	signal k10_needs_bram_8     : bit := '0';
	signal k10_needs_bram_9     : bit := '0';
	signal k10_needs_bram_10     : bit := '0';
	signal k10_needs_bram_11     : bit := '0';
	signal k10_needs_bram_12     : bit := '0';
	signal k10_needs_bram_13     : bit := '0';
	signal k10_needs_bram_14     : bit := '0';
	signal k10_needs_bram_15     : bit := '0';
	signal k11_needs_bram_0     : bit := '0';
	signal k11_needs_bram_1     : bit := '0';
	signal k11_needs_bram_2     : bit := '0';
	signal k11_needs_bram_3     : bit := '0';
	signal k11_needs_bram_4     : bit := '0';
	signal k11_needs_bram_5     : bit := '0';
	signal k11_needs_bram_6     : bit := '0';
	signal k11_needs_bram_7     : bit := '0';
	signal k11_needs_bram_8     : bit := '0';
	signal k11_needs_bram_9     : bit := '0';
	signal k11_needs_bram_10     : bit := '0';
	signal k11_needs_bram_11     : bit := '0';
	signal k11_needs_bram_12     : bit := '0';
	signal k11_needs_bram_13     : bit := '0';
	signal k11_needs_bram_14     : bit := '0';
	signal k11_needs_bram_15     : bit := '0';
	signal k12_needs_bram_0     : bit := '0';
	signal k12_needs_bram_1     : bit := '0';
	signal k12_needs_bram_2     : bit := '0';
	signal k12_needs_bram_3     : bit := '0';
	signal k12_needs_bram_4     : bit := '0';
	signal k12_needs_bram_5     : bit := '0';
	signal k12_needs_bram_6     : bit := '0';
	signal k12_needs_bram_7     : bit := '0';
	signal k12_needs_bram_8     : bit := '0';
	signal k12_needs_bram_9     : bit := '0';
	signal k12_needs_bram_10     : bit := '0';
	signal k12_needs_bram_11     : bit := '0';
	signal k12_needs_bram_12     : bit := '0';
	signal k12_needs_bram_13     : bit := '0';
	signal k12_needs_bram_14     : bit := '0';
	signal k12_needs_bram_15     : bit := '0';
	signal k13_needs_bram_0     : bit := '0';
	signal k13_needs_bram_1     : bit := '0';
	signal k13_needs_bram_2     : bit := '0';
	signal k13_needs_bram_3     : bit := '0';
	signal k13_needs_bram_4     : bit := '0';
	signal k13_needs_bram_5     : bit := '0';
	signal k13_needs_bram_6     : bit := '0';
	signal k13_needs_bram_7     : bit := '0';
	signal k13_needs_bram_8     : bit := '0';
	signal k13_needs_bram_9     : bit := '0';
	signal k13_needs_bram_10     : bit := '0';
	signal k13_needs_bram_11     : bit := '0';
	signal k13_needs_bram_12     : bit := '0';
	signal k13_needs_bram_13     : bit := '0';
	signal k13_needs_bram_14     : bit := '0';
	signal k13_needs_bram_15     : bit := '0';
	signal k14_needs_bram_0     : bit := '0';
	signal k14_needs_bram_1     : bit := '0';
	signal k14_needs_bram_2     : bit := '0';
	signal k14_needs_bram_3     : bit := '0';
	signal k14_needs_bram_4     : bit := '0';
	signal k14_needs_bram_5     : bit := '0';
	signal k14_needs_bram_6     : bit := '0';
	signal k14_needs_bram_7     : bit := '0';
	signal k14_needs_bram_8     : bit := '0';
	signal k14_needs_bram_9     : bit := '0';
	signal k14_needs_bram_10     : bit := '0';
	signal k14_needs_bram_11     : bit := '0';
	signal k14_needs_bram_12     : bit := '0';
	signal k14_needs_bram_13     : bit := '0';
	signal k14_needs_bram_14     : bit := '0';
	signal k14_needs_bram_15     : bit := '0';
	signal k15_needs_bram_0     : bit := '0';
	signal k15_needs_bram_1     : bit := '0';
	signal k15_needs_bram_2     : bit := '0';
	signal k15_needs_bram_3     : bit := '0';
	signal k15_needs_bram_4     : bit := '0';
	signal k15_needs_bram_5     : bit := '0';
	signal k15_needs_bram_6     : bit := '0';
	signal k15_needs_bram_7     : bit := '0';
	signal k15_needs_bram_8     : bit := '0';
	signal k15_needs_bram_9     : bit := '0';
	signal k15_needs_bram_10     : bit := '0';
	signal k15_needs_bram_11     : bit := '0';
	signal k15_needs_bram_12     : bit := '0';
	signal k15_needs_bram_13     : bit := '0';
	signal k15_needs_bram_14     : bit := '0';
	signal k15_needs_bram_15     : bit := '0';
	signal k16_needs_bram_0     : bit := '0';
	signal k16_needs_bram_1     : bit := '0';
	signal k16_needs_bram_2     : bit := '0';
	signal k16_needs_bram_3     : bit := '0';
	signal k16_needs_bram_4     : bit := '0';
	signal k16_needs_bram_5     : bit := '0';
	signal k16_needs_bram_6     : bit := '0';
	signal k16_needs_bram_7     : bit := '0';
	signal k16_needs_bram_8     : bit := '0';
	signal k16_needs_bram_9     : bit := '0';
	signal k16_needs_bram_10     : bit := '0';
	signal k16_needs_bram_11     : bit := '0';
	signal k16_needs_bram_12     : bit := '0';
	signal k16_needs_bram_13     : bit := '0';
	signal k16_needs_bram_14     : bit := '0';
	signal k16_needs_bram_15     : bit := '0';
	signal k17_needs_bram_0     : bit := '0';
	signal k17_needs_bram_1     : bit := '0';
	signal k17_needs_bram_2     : bit := '0';
	signal k17_needs_bram_3     : bit := '0';
	signal k17_needs_bram_4     : bit := '0';
	signal k17_needs_bram_5     : bit := '0';
	signal k17_needs_bram_6     : bit := '0';
	signal k17_needs_bram_7     : bit := '0';
	signal k17_needs_bram_8     : bit := '0';
	signal k17_needs_bram_9     : bit := '0';
	signal k17_needs_bram_10     : bit := '0';
	signal k17_needs_bram_11     : bit := '0';
	signal k17_needs_bram_12     : bit := '0';
	signal k17_needs_bram_13     : bit := '0';
	signal k17_needs_bram_14     : bit := '0';
	signal k17_needs_bram_15     : bit := '0';
	signal k18_needs_bram_0     : bit := '0';
	signal k18_needs_bram_1     : bit := '0';
	signal k18_needs_bram_2     : bit := '0';
	signal k18_needs_bram_3     : bit := '0';
	signal k18_needs_bram_4     : bit := '0';
	signal k18_needs_bram_5     : bit := '0';
	signal k18_needs_bram_6     : bit := '0';
	signal k18_needs_bram_7     : bit := '0';
	signal k18_needs_bram_8     : bit := '0';
	signal k18_needs_bram_9     : bit := '0';
	signal k18_needs_bram_10     : bit := '0';
	signal k18_needs_bram_11     : bit := '0';
	signal k18_needs_bram_12     : bit := '0';
	signal k18_needs_bram_13     : bit := '0';
	signal k18_needs_bram_14     : bit := '0';
	signal k18_needs_bram_15     : bit := '0';
	signal k19_needs_bram_0     : bit := '0';
	signal k19_needs_bram_1     : bit := '0';
	signal k19_needs_bram_2     : bit := '0';
	signal k19_needs_bram_3     : bit := '0';
	signal k19_needs_bram_4     : bit := '0';
	signal k19_needs_bram_5     : bit := '0';
	signal k19_needs_bram_6     : bit := '0';
	signal k19_needs_bram_7     : bit := '0';
	signal k19_needs_bram_8     : bit := '0';
	signal k19_needs_bram_9     : bit := '0';
	signal k19_needs_bram_10     : bit := '0';
	signal k19_needs_bram_11     : bit := '0';
	signal k19_needs_bram_12     : bit := '0';
	signal k19_needs_bram_13     : bit := '0';
	signal k19_needs_bram_14     : bit := '0';
	signal k19_needs_bram_15     : bit := '0';
	signal k20_needs_bram_0     : bit := '0';
	signal k20_needs_bram_1     : bit := '0';
	signal k20_needs_bram_2     : bit := '0';
	signal k20_needs_bram_3     : bit := '0';
	signal k20_needs_bram_4     : bit := '0';
	signal k20_needs_bram_5     : bit := '0';
	signal k20_needs_bram_6     : bit := '0';
	signal k20_needs_bram_7     : bit := '0';
	signal k20_needs_bram_8     : bit := '0';
	signal k20_needs_bram_9     : bit := '0';
	signal k20_needs_bram_10     : bit := '0';
	signal k20_needs_bram_11     : bit := '0';
	signal k20_needs_bram_12     : bit := '0';
	signal k20_needs_bram_13     : bit := '0';
	signal k20_needs_bram_14     : bit := '0';
	signal k20_needs_bram_15     : bit := '0';
	signal k21_needs_bram_0     : bit := '0';
	signal k21_needs_bram_1     : bit := '0';
	signal k21_needs_bram_2     : bit := '0';
	signal k21_needs_bram_3     : bit := '0';
	signal k21_needs_bram_4     : bit := '0';
	signal k21_needs_bram_5     : bit := '0';
	signal k21_needs_bram_6     : bit := '0';
	signal k21_needs_bram_7     : bit := '0';
	signal k21_needs_bram_8     : bit := '0';
	signal k21_needs_bram_9     : bit := '0';
	signal k21_needs_bram_10     : bit := '0';
	signal k21_needs_bram_11     : bit := '0';
	signal k21_needs_bram_12     : bit := '0';
	signal k21_needs_bram_13     : bit := '0';
	signal k21_needs_bram_14     : bit := '0';
	signal k21_needs_bram_15     : bit := '0';
	signal k22_needs_bram_0     : bit := '0';
	signal k22_needs_bram_1     : bit := '0';
	signal k22_needs_bram_2     : bit := '0';
	signal k22_needs_bram_3     : bit := '0';
	signal k22_needs_bram_4     : bit := '0';
	signal k22_needs_bram_5     : bit := '0';
	signal k22_needs_bram_6     : bit := '0';
	signal k22_needs_bram_7     : bit := '0';
	signal k22_needs_bram_8     : bit := '0';
	signal k22_needs_bram_9     : bit := '0';
	signal k22_needs_bram_10     : bit := '0';
	signal k22_needs_bram_11     : bit := '0';
	signal k22_needs_bram_12     : bit := '0';
	signal k22_needs_bram_13     : bit := '0';
	signal k22_needs_bram_14     : bit := '0';
	signal k22_needs_bram_15     : bit := '0';
	signal k23_needs_bram_0     : bit := '0';
	signal k23_needs_bram_1     : bit := '0';
	signal k23_needs_bram_2     : bit := '0';
	signal k23_needs_bram_3     : bit := '0';
	signal k23_needs_bram_4     : bit := '0';
	signal k23_needs_bram_5     : bit := '0';
	signal k23_needs_bram_6     : bit := '0';
	signal k23_needs_bram_7     : bit := '0';
	signal k23_needs_bram_8     : bit := '0';
	signal k23_needs_bram_9     : bit := '0';
	signal k23_needs_bram_10     : bit := '0';
	signal k23_needs_bram_11     : bit := '0';
	signal k23_needs_bram_12     : bit := '0';
	signal k23_needs_bram_13     : bit := '0';
	signal k23_needs_bram_14     : bit := '0';
	signal k23_needs_bram_15     : bit := '0';
	signal k24_needs_bram_0     : bit := '0';
	signal k24_needs_bram_1     : bit := '0';
	signal k24_needs_bram_2     : bit := '0';
	signal k24_needs_bram_3     : bit := '0';
	signal k24_needs_bram_4     : bit := '0';
	signal k24_needs_bram_5     : bit := '0';
	signal k24_needs_bram_6     : bit := '0';
	signal k24_needs_bram_7     : bit := '0';
	signal k24_needs_bram_8     : bit := '0';
	signal k24_needs_bram_9     : bit := '0';
	signal k24_needs_bram_10     : bit := '0';
	signal k24_needs_bram_11     : bit := '0';
	signal k24_needs_bram_12     : bit := '0';
	signal k24_needs_bram_13     : bit := '0';
	signal k24_needs_bram_14     : bit := '0';
	signal k24_needs_bram_15     : bit := '0';
	signal k25_needs_bram_0     : bit := '0';
	signal k25_needs_bram_1     : bit := '0';
	signal k25_needs_bram_2     : bit := '0';
	signal k25_needs_bram_3     : bit := '0';
	signal k25_needs_bram_4     : bit := '0';
	signal k25_needs_bram_5     : bit := '0';
	signal k25_needs_bram_6     : bit := '0';
	signal k25_needs_bram_7     : bit := '0';
	signal k25_needs_bram_8     : bit := '0';
	signal k25_needs_bram_9     : bit := '0';
	signal k25_needs_bram_10     : bit := '0';
	signal k25_needs_bram_11     : bit := '0';
	signal k25_needs_bram_12     : bit := '0';
	signal k25_needs_bram_13     : bit := '0';
	signal k25_needs_bram_14     : bit := '0';
	signal k25_needs_bram_15     : bit := '0';
	signal k26_needs_bram_0     : bit := '0';
	signal k26_needs_bram_1     : bit := '0';
	signal k26_needs_bram_2     : bit := '0';
	signal k26_needs_bram_3     : bit := '0';
	signal k26_needs_bram_4     : bit := '0';
	signal k26_needs_bram_5     : bit := '0';
	signal k26_needs_bram_6     : bit := '0';
	signal k26_needs_bram_7     : bit := '0';
	signal k26_needs_bram_8     : bit := '0';
	signal k26_needs_bram_9     : bit := '0';
	signal k26_needs_bram_10     : bit := '0';
	signal k26_needs_bram_11     : bit := '0';
	signal k26_needs_bram_12     : bit := '0';
	signal k26_needs_bram_13     : bit := '0';
	signal k26_needs_bram_14     : bit := '0';
	signal k26_needs_bram_15     : bit := '0';
	signal k27_needs_bram_0     : bit := '0';
	signal k27_needs_bram_1     : bit := '0';
	signal k27_needs_bram_2     : bit := '0';
	signal k27_needs_bram_3     : bit := '0';
	signal k27_needs_bram_4     : bit := '0';
	signal k27_needs_bram_5     : bit := '0';
	signal k27_needs_bram_6     : bit := '0';
	signal k27_needs_bram_7     : bit := '0';
	signal k27_needs_bram_8     : bit := '0';
	signal k27_needs_bram_9     : bit := '0';
	signal k27_needs_bram_10     : bit := '0';
	signal k27_needs_bram_11     : bit := '0';
	signal k27_needs_bram_12     : bit := '0';
	signal k27_needs_bram_13     : bit := '0';
	signal k27_needs_bram_14     : bit := '0';
	signal k27_needs_bram_15     : bit := '0';
	signal k28_needs_bram_0     : bit := '0';
	signal k28_needs_bram_1     : bit := '0';
	signal k28_needs_bram_2     : bit := '0';
	signal k28_needs_bram_3     : bit := '0';
	signal k28_needs_bram_4     : bit := '0';
	signal k28_needs_bram_5     : bit := '0';
	signal k28_needs_bram_6     : bit := '0';
	signal k28_needs_bram_7     : bit := '0';
	signal k28_needs_bram_8     : bit := '0';
	signal k28_needs_bram_9     : bit := '0';
	signal k28_needs_bram_10     : bit := '0';
	signal k28_needs_bram_11     : bit := '0';
	signal k28_needs_bram_12     : bit := '0';
	signal k28_needs_bram_13     : bit := '0';
	signal k28_needs_bram_14     : bit := '0';
	signal k28_needs_bram_15     : bit := '0';
	signal k29_needs_bram_0     : bit := '0';
	signal k29_needs_bram_1     : bit := '0';
	signal k29_needs_bram_2     : bit := '0';
	signal k29_needs_bram_3     : bit := '0';
	signal k29_needs_bram_4     : bit := '0';
	signal k29_needs_bram_5     : bit := '0';
	signal k29_needs_bram_6     : bit := '0';
	signal k29_needs_bram_7     : bit := '0';
	signal k29_needs_bram_8     : bit := '0';
	signal k29_needs_bram_9     : bit := '0';
	signal k29_needs_bram_10     : bit := '0';
	signal k29_needs_bram_11     : bit := '0';
	signal k29_needs_bram_12     : bit := '0';
	signal k29_needs_bram_13     : bit := '0';
	signal k29_needs_bram_14     : bit := '0';
	signal k29_needs_bram_15     : bit := '0';
	signal k30_needs_bram_0     : bit := '0';
	signal k30_needs_bram_1     : bit := '0';
	signal k30_needs_bram_2     : bit := '0';
	signal k30_needs_bram_3     : bit := '0';
	signal k30_needs_bram_4     : bit := '0';
	signal k30_needs_bram_5     : bit := '0';
	signal k30_needs_bram_6     : bit := '0';
	signal k30_needs_bram_7     : bit := '0';
	signal k30_needs_bram_8     : bit := '0';
	signal k30_needs_bram_9     : bit := '0';
	signal k30_needs_bram_10     : bit := '0';
	signal k30_needs_bram_11     : bit := '0';
	signal k30_needs_bram_12     : bit := '0';
	signal k30_needs_bram_13     : bit := '0';
	signal k30_needs_bram_14     : bit := '0';
	signal k30_needs_bram_15     : bit := '0';
	signal k31_needs_bram_0     : bit := '0';
	signal k31_needs_bram_1     : bit := '0';
	signal k31_needs_bram_2     : bit := '0';
	signal k31_needs_bram_3     : bit := '0';
	signal k31_needs_bram_4     : bit := '0';
	signal k31_needs_bram_5     : bit := '0';
	signal k31_needs_bram_6     : bit := '0';
	signal k31_needs_bram_7     : bit := '0';
	signal k31_needs_bram_8     : bit := '0';
	signal k31_needs_bram_9     : bit := '0';
	signal k31_needs_bram_10     : bit := '0';
	signal k31_needs_bram_11     : bit := '0';
	signal k31_needs_bram_12     : bit := '0';
	signal k31_needs_bram_13     : bit := '0';
	signal k31_needs_bram_14     : bit := '0';
	signal k31_needs_bram_15     : bit := '0';

	signal bram_do             : std_logic_vector(N_PORTS * 32 - 1 downto 0);
	signal bram_di             : std_logic_vector(N_PORTS * 32 - 1 downto 0);
	signal bram_addr           : std_logic_vector(N_PORTS * 9  - 1 downto 0);
	signal bram_we             : std_logic_vector(N_PORTS * 4  - 1 downto 0);
	signal bram_en             : std_logic_vector(N_PORTS * 1  - 1 downto 0);


begin


	bram_en(0) <= '1';
	bram_en(1) <= '1';
	bram_en(2) <= '1';
	bram_en(3) <= '1';
	bram_en(4) <= '1';
	bram_en(5) <= '1';
	bram_en(6) <= '1';
	bram_en(7) <= '1';
	bram_en(8) <= '1';
	bram_en(9) <= '1';
	bram_en(10) <= '1';
	bram_en(11) <= '1';
	bram_en(12) <= '1';
	bram_en(13) <= '1';
	bram_en(14) <= '1';
	bram_en(15) <= '1';
	bram_en(16) <= '1';
	bram_en(17) <= '1';
	bram_en(18) <= '1';
	bram_en(19) <= '1';
	bram_en(20) <= '1';
	bram_en(21) <= '1';
	bram_en(22) <= '1';
	bram_en(23) <= '1';
	bram_en(24) <= '1';
	bram_en(25) <= '1';
	bram_en(26) <= '1';
	bram_en(27) <= '1';
	bram_en(28) <= '1';
	bram_en(29) <= '1';
	bram_en(30) <= '1';
	bram_en(31) <= '1';


	we_0_safe(3) <= WE_0(3) and to_stdulogic(k0_needs_attention);
	we_0_safe(2) <= WE_0(2) and to_stdulogic(k0_needs_attention);
	we_0_safe(1) <= WE_0(1) and to_stdulogic(k0_needs_attention);
	we_0_safe(0) <= WE_0(0) and to_stdulogic(k0_needs_attention);

	we_1_safe(3) <= WE_1(3) and to_stdulogic(k1_needs_attention);
	we_1_safe(2) <= WE_1(2) and to_stdulogic(k1_needs_attention);
	we_1_safe(1) <= WE_1(1) and to_stdulogic(k1_needs_attention);
	we_1_safe(0) <= WE_1(0) and to_stdulogic(k1_needs_attention);

	we_2_safe(3) <= WE_2(3) and to_stdulogic(k2_needs_attention);
	we_2_safe(2) <= WE_2(2) and to_stdulogic(k2_needs_attention);
	we_2_safe(1) <= WE_2(1) and to_stdulogic(k2_needs_attention);
	we_2_safe(0) <= WE_2(0) and to_stdulogic(k2_needs_attention);

	we_3_safe(3) <= WE_3(3) and to_stdulogic(k3_needs_attention);
	we_3_safe(2) <= WE_3(2) and to_stdulogic(k3_needs_attention);
	we_3_safe(1) <= WE_3(1) and to_stdulogic(k3_needs_attention);
	we_3_safe(0) <= WE_3(0) and to_stdulogic(k3_needs_attention);

	we_4_safe(3) <= WE_4(3) and to_stdulogic(k4_needs_attention);
	we_4_safe(2) <= WE_4(2) and to_stdulogic(k4_needs_attention);
	we_4_safe(1) <= WE_4(1) and to_stdulogic(k4_needs_attention);
	we_4_safe(0) <= WE_4(0) and to_stdulogic(k4_needs_attention);

	we_5_safe(3) <= WE_5(3) and to_stdulogic(k5_needs_attention);
	we_5_safe(2) <= WE_5(2) and to_stdulogic(k5_needs_attention);
	we_5_safe(1) <= WE_5(1) and to_stdulogic(k5_needs_attention);
	we_5_safe(0) <= WE_5(0) and to_stdulogic(k5_needs_attention);

	we_6_safe(3) <= WE_6(3) and to_stdulogic(k6_needs_attention);
	we_6_safe(2) <= WE_6(2) and to_stdulogic(k6_needs_attention);
	we_6_safe(1) <= WE_6(1) and to_stdulogic(k6_needs_attention);
	we_6_safe(0) <= WE_6(0) and to_stdulogic(k6_needs_attention);

	we_7_safe(3) <= WE_7(3) and to_stdulogic(k7_needs_attention);
	we_7_safe(2) <= WE_7(2) and to_stdulogic(k7_needs_attention);
	we_7_safe(1) <= WE_7(1) and to_stdulogic(k7_needs_attention);
	we_7_safe(0) <= WE_7(0) and to_stdulogic(k7_needs_attention);

	we_8_safe(3) <= WE_8(3) and to_stdulogic(k8_needs_attention);
	we_8_safe(2) <= WE_8(2) and to_stdulogic(k8_needs_attention);
	we_8_safe(1) <= WE_8(1) and to_stdulogic(k8_needs_attention);
	we_8_safe(0) <= WE_8(0) and to_stdulogic(k8_needs_attention);

	we_9_safe(3) <= WE_9(3) and to_stdulogic(k9_needs_attention);
	we_9_safe(2) <= WE_9(2) and to_stdulogic(k9_needs_attention);
	we_9_safe(1) <= WE_9(1) and to_stdulogic(k9_needs_attention);
	we_9_safe(0) <= WE_9(0) and to_stdulogic(k9_needs_attention);

	we_10_safe(3) <= WE_10(3) and to_stdulogic(k10_needs_attention);
	we_10_safe(2) <= WE_10(2) and to_stdulogic(k10_needs_attention);
	we_10_safe(1) <= WE_10(1) and to_stdulogic(k10_needs_attention);
	we_10_safe(0) <= WE_10(0) and to_stdulogic(k10_needs_attention);

	we_11_safe(3) <= WE_11(3) and to_stdulogic(k11_needs_attention);
	we_11_safe(2) <= WE_11(2) and to_stdulogic(k11_needs_attention);
	we_11_safe(1) <= WE_11(1) and to_stdulogic(k11_needs_attention);
	we_11_safe(0) <= WE_11(0) and to_stdulogic(k11_needs_attention);

	we_12_safe(3) <= WE_12(3) and to_stdulogic(k12_needs_attention);
	we_12_safe(2) <= WE_12(2) and to_stdulogic(k12_needs_attention);
	we_12_safe(1) <= WE_12(1) and to_stdulogic(k12_needs_attention);
	we_12_safe(0) <= WE_12(0) and to_stdulogic(k12_needs_attention);

	we_13_safe(3) <= WE_13(3) and to_stdulogic(k13_needs_attention);
	we_13_safe(2) <= WE_13(2) and to_stdulogic(k13_needs_attention);
	we_13_safe(1) <= WE_13(1) and to_stdulogic(k13_needs_attention);
	we_13_safe(0) <= WE_13(0) and to_stdulogic(k13_needs_attention);

	we_14_safe(3) <= WE_14(3) and to_stdulogic(k14_needs_attention);
	we_14_safe(2) <= WE_14(2) and to_stdulogic(k14_needs_attention);
	we_14_safe(1) <= WE_14(1) and to_stdulogic(k14_needs_attention);
	we_14_safe(0) <= WE_14(0) and to_stdulogic(k14_needs_attention);

	we_15_safe(3) <= WE_15(3) and to_stdulogic(k15_needs_attention);
	we_15_safe(2) <= WE_15(2) and to_stdulogic(k15_needs_attention);
	we_15_safe(1) <= WE_15(1) and to_stdulogic(k15_needs_attention);
	we_15_safe(0) <= WE_15(0) and to_stdulogic(k15_needs_attention);

	we_16_safe(3) <= WE_16(3) and to_stdulogic(k16_needs_attention);
	we_16_safe(2) <= WE_16(2) and to_stdulogic(k16_needs_attention);
	we_16_safe(1) <= WE_16(1) and to_stdulogic(k16_needs_attention);
	we_16_safe(0) <= WE_16(0) and to_stdulogic(k16_needs_attention);

	we_17_safe(3) <= WE_17(3) and to_stdulogic(k17_needs_attention);
	we_17_safe(2) <= WE_17(2) and to_stdulogic(k17_needs_attention);
	we_17_safe(1) <= WE_17(1) and to_stdulogic(k17_needs_attention);
	we_17_safe(0) <= WE_17(0) and to_stdulogic(k17_needs_attention);

	we_18_safe(3) <= WE_18(3) and to_stdulogic(k18_needs_attention);
	we_18_safe(2) <= WE_18(2) and to_stdulogic(k18_needs_attention);
	we_18_safe(1) <= WE_18(1) and to_stdulogic(k18_needs_attention);
	we_18_safe(0) <= WE_18(0) and to_stdulogic(k18_needs_attention);

	we_19_safe(3) <= WE_19(3) and to_stdulogic(k19_needs_attention);
	we_19_safe(2) <= WE_19(2) and to_stdulogic(k19_needs_attention);
	we_19_safe(1) <= WE_19(1) and to_stdulogic(k19_needs_attention);
	we_19_safe(0) <= WE_19(0) and to_stdulogic(k19_needs_attention);

	we_20_safe(3) <= WE_20(3) and to_stdulogic(k20_needs_attention);
	we_20_safe(2) <= WE_20(2) and to_stdulogic(k20_needs_attention);
	we_20_safe(1) <= WE_20(1) and to_stdulogic(k20_needs_attention);
	we_20_safe(0) <= WE_20(0) and to_stdulogic(k20_needs_attention);

	we_21_safe(3) <= WE_21(3) and to_stdulogic(k21_needs_attention);
	we_21_safe(2) <= WE_21(2) and to_stdulogic(k21_needs_attention);
	we_21_safe(1) <= WE_21(1) and to_stdulogic(k21_needs_attention);
	we_21_safe(0) <= WE_21(0) and to_stdulogic(k21_needs_attention);

	we_22_safe(3) <= WE_22(3) and to_stdulogic(k22_needs_attention);
	we_22_safe(2) <= WE_22(2) and to_stdulogic(k22_needs_attention);
	we_22_safe(1) <= WE_22(1) and to_stdulogic(k22_needs_attention);
	we_22_safe(0) <= WE_22(0) and to_stdulogic(k22_needs_attention);

	we_23_safe(3) <= WE_23(3) and to_stdulogic(k23_needs_attention);
	we_23_safe(2) <= WE_23(2) and to_stdulogic(k23_needs_attention);
	we_23_safe(1) <= WE_23(1) and to_stdulogic(k23_needs_attention);
	we_23_safe(0) <= WE_23(0) and to_stdulogic(k23_needs_attention);

	we_24_safe(3) <= WE_24(3) and to_stdulogic(k24_needs_attention);
	we_24_safe(2) <= WE_24(2) and to_stdulogic(k24_needs_attention);
	we_24_safe(1) <= WE_24(1) and to_stdulogic(k24_needs_attention);
	we_24_safe(0) <= WE_24(0) and to_stdulogic(k24_needs_attention);

	we_25_safe(3) <= WE_25(3) and to_stdulogic(k25_needs_attention);
	we_25_safe(2) <= WE_25(2) and to_stdulogic(k25_needs_attention);
	we_25_safe(1) <= WE_25(1) and to_stdulogic(k25_needs_attention);
	we_25_safe(0) <= WE_25(0) and to_stdulogic(k25_needs_attention);

	we_26_safe(3) <= WE_26(3) and to_stdulogic(k26_needs_attention);
	we_26_safe(2) <= WE_26(2) and to_stdulogic(k26_needs_attention);
	we_26_safe(1) <= WE_26(1) and to_stdulogic(k26_needs_attention);
	we_26_safe(0) <= WE_26(0) and to_stdulogic(k26_needs_attention);

	we_27_safe(3) <= WE_27(3) and to_stdulogic(k27_needs_attention);
	we_27_safe(2) <= WE_27(2) and to_stdulogic(k27_needs_attention);
	we_27_safe(1) <= WE_27(1) and to_stdulogic(k27_needs_attention);
	we_27_safe(0) <= WE_27(0) and to_stdulogic(k27_needs_attention);

	we_28_safe(3) <= WE_28(3) and to_stdulogic(k28_needs_attention);
	we_28_safe(2) <= WE_28(2) and to_stdulogic(k28_needs_attention);
	we_28_safe(1) <= WE_28(1) and to_stdulogic(k28_needs_attention);
	we_28_safe(0) <= WE_28(0) and to_stdulogic(k28_needs_attention);

	we_29_safe(3) <= WE_29(3) and to_stdulogic(k29_needs_attention);
	we_29_safe(2) <= WE_29(2) and to_stdulogic(k29_needs_attention);
	we_29_safe(1) <= WE_29(1) and to_stdulogic(k29_needs_attention);
	we_29_safe(0) <= WE_29(0) and to_stdulogic(k29_needs_attention);

	we_30_safe(3) <= WE_30(3) and to_stdulogic(k30_needs_attention);
	we_30_safe(2) <= WE_30(2) and to_stdulogic(k30_needs_attention);
	we_30_safe(1) <= WE_30(1) and to_stdulogic(k30_needs_attention);
	we_30_safe(0) <= WE_30(0) and to_stdulogic(k30_needs_attention);

	we_31_safe(3) <= WE_31(3) and to_stdulogic(k31_needs_attention);
	we_31_safe(2) <= WE_31(2) and to_stdulogic(k31_needs_attention);
	we_31_safe(1) <= WE_31(1) and to_stdulogic(k31_needs_attention);
	we_31_safe(0) <= WE_31(0) and to_stdulogic(k31_needs_attention);


	RDY_0 <= to_stdulogic(k0_being_served);
	RDY_1 <= to_stdulogic(k1_being_served);
	RDY_2 <= to_stdulogic(k2_being_served);
	RDY_3 <= to_stdulogic(k3_being_served);
	RDY_4 <= to_stdulogic(k4_being_served);
	RDY_5 <= to_stdulogic(k5_being_served);
	RDY_6 <= to_stdulogic(k6_being_served);
	RDY_7 <= to_stdulogic(k7_being_served);
	RDY_8 <= to_stdulogic(k8_being_served);
	RDY_9 <= to_stdulogic(k9_being_served);
	RDY_10 <= to_stdulogic(k10_being_served);
	RDY_11 <= to_stdulogic(k11_being_served);
	RDY_12 <= to_stdulogic(k12_being_served);
	RDY_13 <= to_stdulogic(k13_being_served);
	RDY_14 <= to_stdulogic(k14_being_served);
	RDY_15 <= to_stdulogic(k15_being_served);
	RDY_16 <= to_stdulogic(k16_being_served);
	RDY_17 <= to_stdulogic(k17_being_served);
	RDY_18 <= to_stdulogic(k18_being_served);
	RDY_19 <= to_stdulogic(k19_being_served);
	RDY_20 <= to_stdulogic(k20_being_served);
	RDY_21 <= to_stdulogic(k21_being_served);
	RDY_22 <= to_stdulogic(k22_being_served);
	RDY_23 <= to_stdulogic(k23_being_served);
	RDY_24 <= to_stdulogic(k24_being_served);
	RDY_25 <= to_stdulogic(k25_being_served);
	RDY_26 <= to_stdulogic(k26_being_served);
	RDY_27 <= to_stdulogic(k27_being_served);
	RDY_28 <= to_stdulogic(k28_being_served);
	RDY_29 <= to_stdulogic(k29_being_served);
	RDY_30 <= to_stdulogic(k30_being_served);
	RDY_31 <= to_stdulogic(k31_being_served);


	k0_needs_attention <= to_bit(REQ_0);

	k1_needs_attention <= to_bit(REQ_1) and (not (addr_0_eq_addr_1 and k0_needs_attention));

	k2_needs_attention <= to_bit(REQ_2) and (not (addr_0_eq_addr_2 and k0_needs_attention)) and (not (addr_1_eq_addr_2 and k1_needs_attention));

	k3_needs_attention <= to_bit(REQ_3) and (not (addr_0_eq_addr_3 and k0_needs_attention)) and (not (addr_1_eq_addr_3 and k1_needs_attention)) and (not (addr_2_eq_addr_3 and k2_needs_attention));

	k4_needs_attention <= to_bit(REQ_4) and (not (addr_0_eq_addr_4 and k0_needs_attention)) and (not (addr_1_eq_addr_4 and k1_needs_attention)) and (not (addr_2_eq_addr_4 and k2_needs_attention)) and (not (addr_3_eq_addr_4 and k3_needs_attention));

	k5_needs_attention <= to_bit(REQ_5) and (not (addr_0_eq_addr_5 and k0_needs_attention)) and (not (addr_1_eq_addr_5 and k1_needs_attention)) and (not (addr_2_eq_addr_5 and k2_needs_attention)) and (not (addr_3_eq_addr_5 and k3_needs_attention)) and (not (addr_4_eq_addr_5 and k4_needs_attention));

	k6_needs_attention <= to_bit(REQ_6) and (not (addr_0_eq_addr_6 and k0_needs_attention)) and (not (addr_1_eq_addr_6 and k1_needs_attention)) and (not (addr_2_eq_addr_6 and k2_needs_attention)) and (not (addr_3_eq_addr_6 and k3_needs_attention)) and (not (addr_4_eq_addr_6 and k4_needs_attention)) and (not (addr_5_eq_addr_6 and k5_needs_attention));

	k7_needs_attention <= to_bit(REQ_7) and (not (addr_0_eq_addr_7 and k0_needs_attention)) and (not (addr_1_eq_addr_7 and k1_needs_attention)) and (not (addr_2_eq_addr_7 and k2_needs_attention)) and (not (addr_3_eq_addr_7 and k3_needs_attention)) and (not (addr_4_eq_addr_7 and k4_needs_attention)) and (not (addr_5_eq_addr_7 and k5_needs_attention)) and (not (addr_6_eq_addr_7 and k6_needs_attention));

	k8_needs_attention <= to_bit(REQ_8) and (not (addr_0_eq_addr_8 and k0_needs_attention)) and (not (addr_1_eq_addr_8 and k1_needs_attention)) and (not (addr_2_eq_addr_8 and k2_needs_attention)) and (not (addr_3_eq_addr_8 and k3_needs_attention)) and (not (addr_4_eq_addr_8 and k4_needs_attention)) and (not (addr_5_eq_addr_8 and k5_needs_attention)) and (not (addr_6_eq_addr_8 and k6_needs_attention)) and (not (addr_7_eq_addr_8 and k7_needs_attention));

	k9_needs_attention <= to_bit(REQ_9) and (not (addr_0_eq_addr_9 and k0_needs_attention)) and (not (addr_1_eq_addr_9 and k1_needs_attention)) and (not (addr_2_eq_addr_9 and k2_needs_attention)) and (not (addr_3_eq_addr_9 and k3_needs_attention)) and (not (addr_4_eq_addr_9 and k4_needs_attention)) and (not (addr_5_eq_addr_9 and k5_needs_attention)) and (not (addr_6_eq_addr_9 and k6_needs_attention)) and (not (addr_7_eq_addr_9 and k7_needs_attention)) and (not (addr_8_eq_addr_9 and k8_needs_attention));

	k10_needs_attention <= to_bit(REQ_10) and (not (addr_0_eq_addr_10 and k0_needs_attention)) and (not (addr_1_eq_addr_10 and k1_needs_attention)) and (not (addr_2_eq_addr_10 and k2_needs_attention)) and (not (addr_3_eq_addr_10 and k3_needs_attention)) and (not (addr_4_eq_addr_10 and k4_needs_attention)) and (not (addr_5_eq_addr_10 and k5_needs_attention)) and (not (addr_6_eq_addr_10 and k6_needs_attention)) and (not (addr_7_eq_addr_10 and k7_needs_attention)) and (not (addr_8_eq_addr_10 and k8_needs_attention)) and (not (addr_9_eq_addr_10 and k9_needs_attention));

	k11_needs_attention <= to_bit(REQ_11) and (not (addr_0_eq_addr_11 and k0_needs_attention)) and (not (addr_1_eq_addr_11 and k1_needs_attention)) and (not (addr_2_eq_addr_11 and k2_needs_attention)) and (not (addr_3_eq_addr_11 and k3_needs_attention)) and (not (addr_4_eq_addr_11 and k4_needs_attention)) and (not (addr_5_eq_addr_11 and k5_needs_attention)) and (not (addr_6_eq_addr_11 and k6_needs_attention)) and (not (addr_7_eq_addr_11 and k7_needs_attention)) and (not (addr_8_eq_addr_11 and k8_needs_attention)) and (not (addr_9_eq_addr_11 and k9_needs_attention)) and (not (addr_10_eq_addr_11 and k10_needs_attention));

	k12_needs_attention <= to_bit(REQ_12) and (not (addr_0_eq_addr_12 and k0_needs_attention)) and (not (addr_1_eq_addr_12 and k1_needs_attention)) and (not (addr_2_eq_addr_12 and k2_needs_attention)) and (not (addr_3_eq_addr_12 and k3_needs_attention)) and (not (addr_4_eq_addr_12 and k4_needs_attention)) and (not (addr_5_eq_addr_12 and k5_needs_attention)) and (not (addr_6_eq_addr_12 and k6_needs_attention)) and (not (addr_7_eq_addr_12 and k7_needs_attention)) and (not (addr_8_eq_addr_12 and k8_needs_attention)) and (not (addr_9_eq_addr_12 and k9_needs_attention)) and (not (addr_10_eq_addr_12 and k10_needs_attention)) and (not (addr_11_eq_addr_12 and k11_needs_attention));

	k13_needs_attention <= to_bit(REQ_13) and (not (addr_0_eq_addr_13 and k0_needs_attention)) and (not (addr_1_eq_addr_13 and k1_needs_attention)) and (not (addr_2_eq_addr_13 and k2_needs_attention)) and (not (addr_3_eq_addr_13 and k3_needs_attention)) and (not (addr_4_eq_addr_13 and k4_needs_attention)) and (not (addr_5_eq_addr_13 and k5_needs_attention)) and (not (addr_6_eq_addr_13 and k6_needs_attention)) and (not (addr_7_eq_addr_13 and k7_needs_attention)) and (not (addr_8_eq_addr_13 and k8_needs_attention)) and (not (addr_9_eq_addr_13 and k9_needs_attention)) and (not (addr_10_eq_addr_13 and k10_needs_attention)) and (not (addr_11_eq_addr_13 and k11_needs_attention)) and (not (addr_12_eq_addr_13 and k12_needs_attention));

	k14_needs_attention <= to_bit(REQ_14) and (not (addr_0_eq_addr_14 and k0_needs_attention)) and (not (addr_1_eq_addr_14 and k1_needs_attention)) and (not (addr_2_eq_addr_14 and k2_needs_attention)) and (not (addr_3_eq_addr_14 and k3_needs_attention)) and (not (addr_4_eq_addr_14 and k4_needs_attention)) and (not (addr_5_eq_addr_14 and k5_needs_attention)) and (not (addr_6_eq_addr_14 and k6_needs_attention)) and (not (addr_7_eq_addr_14 and k7_needs_attention)) and (not (addr_8_eq_addr_14 and k8_needs_attention)) and (not (addr_9_eq_addr_14 and k9_needs_attention)) and (not (addr_10_eq_addr_14 and k10_needs_attention)) and (not (addr_11_eq_addr_14 and k11_needs_attention)) and (not (addr_12_eq_addr_14 and k12_needs_attention)) and (not (addr_13_eq_addr_14 and k13_needs_attention));

	k15_needs_attention <= to_bit(REQ_15) and (not (addr_0_eq_addr_15 and k0_needs_attention)) and (not (addr_1_eq_addr_15 and k1_needs_attention)) and (not (addr_2_eq_addr_15 and k2_needs_attention)) and (not (addr_3_eq_addr_15 and k3_needs_attention)) and (not (addr_4_eq_addr_15 and k4_needs_attention)) and (not (addr_5_eq_addr_15 and k5_needs_attention)) and (not (addr_6_eq_addr_15 and k6_needs_attention)) and (not (addr_7_eq_addr_15 and k7_needs_attention)) and (not (addr_8_eq_addr_15 and k8_needs_attention)) and (not (addr_9_eq_addr_15 and k9_needs_attention)) and (not (addr_10_eq_addr_15 and k10_needs_attention)) and (not (addr_11_eq_addr_15 and k11_needs_attention)) and (not (addr_12_eq_addr_15 and k12_needs_attention)) and (not (addr_13_eq_addr_15 and k13_needs_attention)) and (not (addr_14_eq_addr_15 and k14_needs_attention));

	k16_needs_attention <= to_bit(REQ_16) and (not (addr_0_eq_addr_16 and k0_needs_attention)) and (not (addr_1_eq_addr_16 and k1_needs_attention)) and (not (addr_2_eq_addr_16 and k2_needs_attention)) and (not (addr_3_eq_addr_16 and k3_needs_attention)) and (not (addr_4_eq_addr_16 and k4_needs_attention)) and (not (addr_5_eq_addr_16 and k5_needs_attention)) and (not (addr_6_eq_addr_16 and k6_needs_attention)) and (not (addr_7_eq_addr_16 and k7_needs_attention)) and (not (addr_8_eq_addr_16 and k8_needs_attention)) and (not (addr_9_eq_addr_16 and k9_needs_attention)) and (not (addr_10_eq_addr_16 and k10_needs_attention)) and (not (addr_11_eq_addr_16 and k11_needs_attention)) and (not (addr_12_eq_addr_16 and k12_needs_attention)) and (not (addr_13_eq_addr_16 and k13_needs_attention)) and (not (addr_14_eq_addr_16 and k14_needs_attention)) and (not (addr_15_eq_addr_16 and k15_needs_attention));

	k17_needs_attention <= to_bit(REQ_17) and (not (addr_0_eq_addr_17 and k0_needs_attention)) and (not (addr_1_eq_addr_17 and k1_needs_attention)) and (not (addr_2_eq_addr_17 and k2_needs_attention)) and (not (addr_3_eq_addr_17 and k3_needs_attention)) and (not (addr_4_eq_addr_17 and k4_needs_attention)) and (not (addr_5_eq_addr_17 and k5_needs_attention)) and (not (addr_6_eq_addr_17 and k6_needs_attention)) and (not (addr_7_eq_addr_17 and k7_needs_attention)) and (not (addr_8_eq_addr_17 and k8_needs_attention)) and (not (addr_9_eq_addr_17 and k9_needs_attention)) and (not (addr_10_eq_addr_17 and k10_needs_attention)) and (not (addr_11_eq_addr_17 and k11_needs_attention)) and (not (addr_12_eq_addr_17 and k12_needs_attention)) and (not (addr_13_eq_addr_17 and k13_needs_attention)) and (not (addr_14_eq_addr_17 and k14_needs_attention)) and (not (addr_15_eq_addr_17 and k15_needs_attention)) and (not (addr_16_eq_addr_17 and k16_needs_attention));

	k18_needs_attention <= to_bit(REQ_18) and (not (addr_0_eq_addr_18 and k0_needs_attention)) and (not (addr_1_eq_addr_18 and k1_needs_attention)) and (not (addr_2_eq_addr_18 and k2_needs_attention)) and (not (addr_3_eq_addr_18 and k3_needs_attention)) and (not (addr_4_eq_addr_18 and k4_needs_attention)) and (not (addr_5_eq_addr_18 and k5_needs_attention)) and (not (addr_6_eq_addr_18 and k6_needs_attention)) and (not (addr_7_eq_addr_18 and k7_needs_attention)) and (not (addr_8_eq_addr_18 and k8_needs_attention)) and (not (addr_9_eq_addr_18 and k9_needs_attention)) and (not (addr_10_eq_addr_18 and k10_needs_attention)) and (not (addr_11_eq_addr_18 and k11_needs_attention)) and (not (addr_12_eq_addr_18 and k12_needs_attention)) and (not (addr_13_eq_addr_18 and k13_needs_attention)) and (not (addr_14_eq_addr_18 and k14_needs_attention)) and (not (addr_15_eq_addr_18 and k15_needs_attention)) and (not (addr_16_eq_addr_18 and k16_needs_attention)) and (not (addr_17_eq_addr_18 and k17_needs_attention));

	k19_needs_attention <= to_bit(REQ_19) and (not (addr_0_eq_addr_19 and k0_needs_attention)) and (not (addr_1_eq_addr_19 and k1_needs_attention)) and (not (addr_2_eq_addr_19 and k2_needs_attention)) and (not (addr_3_eq_addr_19 and k3_needs_attention)) and (not (addr_4_eq_addr_19 and k4_needs_attention)) and (not (addr_5_eq_addr_19 and k5_needs_attention)) and (not (addr_6_eq_addr_19 and k6_needs_attention)) and (not (addr_7_eq_addr_19 and k7_needs_attention)) and (not (addr_8_eq_addr_19 and k8_needs_attention)) and (not (addr_9_eq_addr_19 and k9_needs_attention)) and (not (addr_10_eq_addr_19 and k10_needs_attention)) and (not (addr_11_eq_addr_19 and k11_needs_attention)) and (not (addr_12_eq_addr_19 and k12_needs_attention)) and (not (addr_13_eq_addr_19 and k13_needs_attention)) and (not (addr_14_eq_addr_19 and k14_needs_attention)) and (not (addr_15_eq_addr_19 and k15_needs_attention)) and (not (addr_16_eq_addr_19 and k16_needs_attention)) and (not (addr_17_eq_addr_19 and k17_needs_attention)) and (not (addr_18_eq_addr_19 and k18_needs_attention));

	k20_needs_attention <= to_bit(REQ_20) and (not (addr_0_eq_addr_20 and k0_needs_attention)) and (not (addr_1_eq_addr_20 and k1_needs_attention)) and (not (addr_2_eq_addr_20 and k2_needs_attention)) and (not (addr_3_eq_addr_20 and k3_needs_attention)) and (not (addr_4_eq_addr_20 and k4_needs_attention)) and (not (addr_5_eq_addr_20 and k5_needs_attention)) and (not (addr_6_eq_addr_20 and k6_needs_attention)) and (not (addr_7_eq_addr_20 and k7_needs_attention)) and (not (addr_8_eq_addr_20 and k8_needs_attention)) and (not (addr_9_eq_addr_20 and k9_needs_attention)) and (not (addr_10_eq_addr_20 and k10_needs_attention)) and (not (addr_11_eq_addr_20 and k11_needs_attention)) and (not (addr_12_eq_addr_20 and k12_needs_attention)) and (not (addr_13_eq_addr_20 and k13_needs_attention)) and (not (addr_14_eq_addr_20 and k14_needs_attention)) and (not (addr_15_eq_addr_20 and k15_needs_attention)) and (not (addr_16_eq_addr_20 and k16_needs_attention)) and (not (addr_17_eq_addr_20 and k17_needs_attention)) and (not (addr_18_eq_addr_20 and k18_needs_attention)) and (not (addr_19_eq_addr_20 and k19_needs_attention));

	k21_needs_attention <= to_bit(REQ_21) and (not (addr_0_eq_addr_21 and k0_needs_attention)) and (not (addr_1_eq_addr_21 and k1_needs_attention)) and (not (addr_2_eq_addr_21 and k2_needs_attention)) and (not (addr_3_eq_addr_21 and k3_needs_attention)) and (not (addr_4_eq_addr_21 and k4_needs_attention)) and (not (addr_5_eq_addr_21 and k5_needs_attention)) and (not (addr_6_eq_addr_21 and k6_needs_attention)) and (not (addr_7_eq_addr_21 and k7_needs_attention)) and (not (addr_8_eq_addr_21 and k8_needs_attention)) and (not (addr_9_eq_addr_21 and k9_needs_attention)) and (not (addr_10_eq_addr_21 and k10_needs_attention)) and (not (addr_11_eq_addr_21 and k11_needs_attention)) and (not (addr_12_eq_addr_21 and k12_needs_attention)) and (not (addr_13_eq_addr_21 and k13_needs_attention)) and (not (addr_14_eq_addr_21 and k14_needs_attention)) and (not (addr_15_eq_addr_21 and k15_needs_attention)) and (not (addr_16_eq_addr_21 and k16_needs_attention)) and (not (addr_17_eq_addr_21 and k17_needs_attention)) and (not (addr_18_eq_addr_21 and k18_needs_attention)) and (not (addr_19_eq_addr_21 and k19_needs_attention)) and (not (addr_20_eq_addr_21 and k20_needs_attention));

	k22_needs_attention <= to_bit(REQ_22) and (not (addr_0_eq_addr_22 and k0_needs_attention)) and (not (addr_1_eq_addr_22 and k1_needs_attention)) and (not (addr_2_eq_addr_22 and k2_needs_attention)) and (not (addr_3_eq_addr_22 and k3_needs_attention)) and (not (addr_4_eq_addr_22 and k4_needs_attention)) and (not (addr_5_eq_addr_22 and k5_needs_attention)) and (not (addr_6_eq_addr_22 and k6_needs_attention)) and (not (addr_7_eq_addr_22 and k7_needs_attention)) and (not (addr_8_eq_addr_22 and k8_needs_attention)) and (not (addr_9_eq_addr_22 and k9_needs_attention)) and (not (addr_10_eq_addr_22 and k10_needs_attention)) and (not (addr_11_eq_addr_22 and k11_needs_attention)) and (not (addr_12_eq_addr_22 and k12_needs_attention)) and (not (addr_13_eq_addr_22 and k13_needs_attention)) and (not (addr_14_eq_addr_22 and k14_needs_attention)) and (not (addr_15_eq_addr_22 and k15_needs_attention)) and (not (addr_16_eq_addr_22 and k16_needs_attention)) and (not (addr_17_eq_addr_22 and k17_needs_attention)) and (not (addr_18_eq_addr_22 and k18_needs_attention)) and (not (addr_19_eq_addr_22 and k19_needs_attention)) and (not (addr_20_eq_addr_22 and k20_needs_attention)) and (not (addr_21_eq_addr_22 and k21_needs_attention));

	k23_needs_attention <= to_bit(REQ_23) and (not (addr_0_eq_addr_23 and k0_needs_attention)) and (not (addr_1_eq_addr_23 and k1_needs_attention)) and (not (addr_2_eq_addr_23 and k2_needs_attention)) and (not (addr_3_eq_addr_23 and k3_needs_attention)) and (not (addr_4_eq_addr_23 and k4_needs_attention)) and (not (addr_5_eq_addr_23 and k5_needs_attention)) and (not (addr_6_eq_addr_23 and k6_needs_attention)) and (not (addr_7_eq_addr_23 and k7_needs_attention)) and (not (addr_8_eq_addr_23 and k8_needs_attention)) and (not (addr_9_eq_addr_23 and k9_needs_attention)) and (not (addr_10_eq_addr_23 and k10_needs_attention)) and (not (addr_11_eq_addr_23 and k11_needs_attention)) and (not (addr_12_eq_addr_23 and k12_needs_attention)) and (not (addr_13_eq_addr_23 and k13_needs_attention)) and (not (addr_14_eq_addr_23 and k14_needs_attention)) and (not (addr_15_eq_addr_23 and k15_needs_attention)) and (not (addr_16_eq_addr_23 and k16_needs_attention)) and (not (addr_17_eq_addr_23 and k17_needs_attention)) and (not (addr_18_eq_addr_23 and k18_needs_attention)) and (not (addr_19_eq_addr_23 and k19_needs_attention)) and (not (addr_20_eq_addr_23 and k20_needs_attention)) and (not (addr_21_eq_addr_23 and k21_needs_attention)) and (not (addr_22_eq_addr_23 and k22_needs_attention));

	k24_needs_attention <= to_bit(REQ_24) and (not (addr_0_eq_addr_24 and k0_needs_attention)) and (not (addr_1_eq_addr_24 and k1_needs_attention)) and (not (addr_2_eq_addr_24 and k2_needs_attention)) and (not (addr_3_eq_addr_24 and k3_needs_attention)) and (not (addr_4_eq_addr_24 and k4_needs_attention)) and (not (addr_5_eq_addr_24 and k5_needs_attention)) and (not (addr_6_eq_addr_24 and k6_needs_attention)) and (not (addr_7_eq_addr_24 and k7_needs_attention)) and (not (addr_8_eq_addr_24 and k8_needs_attention)) and (not (addr_9_eq_addr_24 and k9_needs_attention)) and (not (addr_10_eq_addr_24 and k10_needs_attention)) and (not (addr_11_eq_addr_24 and k11_needs_attention)) and (not (addr_12_eq_addr_24 and k12_needs_attention)) and (not (addr_13_eq_addr_24 and k13_needs_attention)) and (not (addr_14_eq_addr_24 and k14_needs_attention)) and (not (addr_15_eq_addr_24 and k15_needs_attention)) and (not (addr_16_eq_addr_24 and k16_needs_attention)) and (not (addr_17_eq_addr_24 and k17_needs_attention)) and (not (addr_18_eq_addr_24 and k18_needs_attention)) and (not (addr_19_eq_addr_24 and k19_needs_attention)) and (not (addr_20_eq_addr_24 and k20_needs_attention)) and (not (addr_21_eq_addr_24 and k21_needs_attention)) and (not (addr_22_eq_addr_24 and k22_needs_attention)) and (not (addr_23_eq_addr_24 and k23_needs_attention));

	k25_needs_attention <= to_bit(REQ_25) and (not (addr_0_eq_addr_25 and k0_needs_attention)) and (not (addr_1_eq_addr_25 and k1_needs_attention)) and (not (addr_2_eq_addr_25 and k2_needs_attention)) and (not (addr_3_eq_addr_25 and k3_needs_attention)) and (not (addr_4_eq_addr_25 and k4_needs_attention)) and (not (addr_5_eq_addr_25 and k5_needs_attention)) and (not (addr_6_eq_addr_25 and k6_needs_attention)) and (not (addr_7_eq_addr_25 and k7_needs_attention)) and (not (addr_8_eq_addr_25 and k8_needs_attention)) and (not (addr_9_eq_addr_25 and k9_needs_attention)) and (not (addr_10_eq_addr_25 and k10_needs_attention)) and (not (addr_11_eq_addr_25 and k11_needs_attention)) and (not (addr_12_eq_addr_25 and k12_needs_attention)) and (not (addr_13_eq_addr_25 and k13_needs_attention)) and (not (addr_14_eq_addr_25 and k14_needs_attention)) and (not (addr_15_eq_addr_25 and k15_needs_attention)) and (not (addr_16_eq_addr_25 and k16_needs_attention)) and (not (addr_17_eq_addr_25 and k17_needs_attention)) and (not (addr_18_eq_addr_25 and k18_needs_attention)) and (not (addr_19_eq_addr_25 and k19_needs_attention)) and (not (addr_20_eq_addr_25 and k20_needs_attention)) and (not (addr_21_eq_addr_25 and k21_needs_attention)) and (not (addr_22_eq_addr_25 and k22_needs_attention)) and (not (addr_23_eq_addr_25 and k23_needs_attention)) and (not (addr_24_eq_addr_25 and k24_needs_attention));

	k26_needs_attention <= to_bit(REQ_26) and (not (addr_0_eq_addr_26 and k0_needs_attention)) and (not (addr_1_eq_addr_26 and k1_needs_attention)) and (not (addr_2_eq_addr_26 and k2_needs_attention)) and (not (addr_3_eq_addr_26 and k3_needs_attention)) and (not (addr_4_eq_addr_26 and k4_needs_attention)) and (not (addr_5_eq_addr_26 and k5_needs_attention)) and (not (addr_6_eq_addr_26 and k6_needs_attention)) and (not (addr_7_eq_addr_26 and k7_needs_attention)) and (not (addr_8_eq_addr_26 and k8_needs_attention)) and (not (addr_9_eq_addr_26 and k9_needs_attention)) and (not (addr_10_eq_addr_26 and k10_needs_attention)) and (not (addr_11_eq_addr_26 and k11_needs_attention)) and (not (addr_12_eq_addr_26 and k12_needs_attention)) and (not (addr_13_eq_addr_26 and k13_needs_attention)) and (not (addr_14_eq_addr_26 and k14_needs_attention)) and (not (addr_15_eq_addr_26 and k15_needs_attention)) and (not (addr_16_eq_addr_26 and k16_needs_attention)) and (not (addr_17_eq_addr_26 and k17_needs_attention)) and (not (addr_18_eq_addr_26 and k18_needs_attention)) and (not (addr_19_eq_addr_26 and k19_needs_attention)) and (not (addr_20_eq_addr_26 and k20_needs_attention)) and (not (addr_21_eq_addr_26 and k21_needs_attention)) and (not (addr_22_eq_addr_26 and k22_needs_attention)) and (not (addr_23_eq_addr_26 and k23_needs_attention)) and (not (addr_24_eq_addr_26 and k24_needs_attention)) and (not (addr_25_eq_addr_26 and k25_needs_attention));

	k27_needs_attention <= to_bit(REQ_27) and (not (addr_0_eq_addr_27 and k0_needs_attention)) and (not (addr_1_eq_addr_27 and k1_needs_attention)) and (not (addr_2_eq_addr_27 and k2_needs_attention)) and (not (addr_3_eq_addr_27 and k3_needs_attention)) and (not (addr_4_eq_addr_27 and k4_needs_attention)) and (not (addr_5_eq_addr_27 and k5_needs_attention)) and (not (addr_6_eq_addr_27 and k6_needs_attention)) and (not (addr_7_eq_addr_27 and k7_needs_attention)) and (not (addr_8_eq_addr_27 and k8_needs_attention)) and (not (addr_9_eq_addr_27 and k9_needs_attention)) and (not (addr_10_eq_addr_27 and k10_needs_attention)) and (not (addr_11_eq_addr_27 and k11_needs_attention)) and (not (addr_12_eq_addr_27 and k12_needs_attention)) and (not (addr_13_eq_addr_27 and k13_needs_attention)) and (not (addr_14_eq_addr_27 and k14_needs_attention)) and (not (addr_15_eq_addr_27 and k15_needs_attention)) and (not (addr_16_eq_addr_27 and k16_needs_attention)) and (not (addr_17_eq_addr_27 and k17_needs_attention)) and (not (addr_18_eq_addr_27 and k18_needs_attention)) and (not (addr_19_eq_addr_27 and k19_needs_attention)) and (not (addr_20_eq_addr_27 and k20_needs_attention)) and (not (addr_21_eq_addr_27 and k21_needs_attention)) and (not (addr_22_eq_addr_27 and k22_needs_attention)) and (not (addr_23_eq_addr_27 and k23_needs_attention)) and (not (addr_24_eq_addr_27 and k24_needs_attention)) and (not (addr_25_eq_addr_27 and k25_needs_attention)) and (not (addr_26_eq_addr_27 and k26_needs_attention));

	k28_needs_attention <= to_bit(REQ_28) and (not (addr_0_eq_addr_28 and k0_needs_attention)) and (not (addr_1_eq_addr_28 and k1_needs_attention)) and (not (addr_2_eq_addr_28 and k2_needs_attention)) and (not (addr_3_eq_addr_28 and k3_needs_attention)) and (not (addr_4_eq_addr_28 and k4_needs_attention)) and (not (addr_5_eq_addr_28 and k5_needs_attention)) and (not (addr_6_eq_addr_28 and k6_needs_attention)) and (not (addr_7_eq_addr_28 and k7_needs_attention)) and (not (addr_8_eq_addr_28 and k8_needs_attention)) and (not (addr_9_eq_addr_28 and k9_needs_attention)) and (not (addr_10_eq_addr_28 and k10_needs_attention)) and (not (addr_11_eq_addr_28 and k11_needs_attention)) and (not (addr_12_eq_addr_28 and k12_needs_attention)) and (not (addr_13_eq_addr_28 and k13_needs_attention)) and (not (addr_14_eq_addr_28 and k14_needs_attention)) and (not (addr_15_eq_addr_28 and k15_needs_attention)) and (not (addr_16_eq_addr_28 and k16_needs_attention)) and (not (addr_17_eq_addr_28 and k17_needs_attention)) and (not (addr_18_eq_addr_28 and k18_needs_attention)) and (not (addr_19_eq_addr_28 and k19_needs_attention)) and (not (addr_20_eq_addr_28 and k20_needs_attention)) and (not (addr_21_eq_addr_28 and k21_needs_attention)) and (not (addr_22_eq_addr_28 and k22_needs_attention)) and (not (addr_23_eq_addr_28 and k23_needs_attention)) and (not (addr_24_eq_addr_28 and k24_needs_attention)) and (not (addr_25_eq_addr_28 and k25_needs_attention)) and (not (addr_26_eq_addr_28 and k26_needs_attention)) and (not (addr_27_eq_addr_28 and k27_needs_attention));

	k29_needs_attention <= to_bit(REQ_29) and (not (addr_0_eq_addr_29 and k0_needs_attention)) and (not (addr_1_eq_addr_29 and k1_needs_attention)) and (not (addr_2_eq_addr_29 and k2_needs_attention)) and (not (addr_3_eq_addr_29 and k3_needs_attention)) and (not (addr_4_eq_addr_29 and k4_needs_attention)) and (not (addr_5_eq_addr_29 and k5_needs_attention)) and (not (addr_6_eq_addr_29 and k6_needs_attention)) and (not (addr_7_eq_addr_29 and k7_needs_attention)) and (not (addr_8_eq_addr_29 and k8_needs_attention)) and (not (addr_9_eq_addr_29 and k9_needs_attention)) and (not (addr_10_eq_addr_29 and k10_needs_attention)) and (not (addr_11_eq_addr_29 and k11_needs_attention)) and (not (addr_12_eq_addr_29 and k12_needs_attention)) and (not (addr_13_eq_addr_29 and k13_needs_attention)) and (not (addr_14_eq_addr_29 and k14_needs_attention)) and (not (addr_15_eq_addr_29 and k15_needs_attention)) and (not (addr_16_eq_addr_29 and k16_needs_attention)) and (not (addr_17_eq_addr_29 and k17_needs_attention)) and (not (addr_18_eq_addr_29 and k18_needs_attention)) and (not (addr_19_eq_addr_29 and k19_needs_attention)) and (not (addr_20_eq_addr_29 and k20_needs_attention)) and (not (addr_21_eq_addr_29 and k21_needs_attention)) and (not (addr_22_eq_addr_29 and k22_needs_attention)) and (not (addr_23_eq_addr_29 and k23_needs_attention)) and (not (addr_24_eq_addr_29 and k24_needs_attention)) and (not (addr_25_eq_addr_29 and k25_needs_attention)) and (not (addr_26_eq_addr_29 and k26_needs_attention)) and (not (addr_27_eq_addr_29 and k27_needs_attention)) and (not (addr_28_eq_addr_29 and k28_needs_attention));

	k30_needs_attention <= to_bit(REQ_30) and (not (addr_0_eq_addr_30 and k0_needs_attention)) and (not (addr_1_eq_addr_30 and k1_needs_attention)) and (not (addr_2_eq_addr_30 and k2_needs_attention)) and (not (addr_3_eq_addr_30 and k3_needs_attention)) and (not (addr_4_eq_addr_30 and k4_needs_attention)) and (not (addr_5_eq_addr_30 and k5_needs_attention)) and (not (addr_6_eq_addr_30 and k6_needs_attention)) and (not (addr_7_eq_addr_30 and k7_needs_attention)) and (not (addr_8_eq_addr_30 and k8_needs_attention)) and (not (addr_9_eq_addr_30 and k9_needs_attention)) and (not (addr_10_eq_addr_30 and k10_needs_attention)) and (not (addr_11_eq_addr_30 and k11_needs_attention)) and (not (addr_12_eq_addr_30 and k12_needs_attention)) and (not (addr_13_eq_addr_30 and k13_needs_attention)) and (not (addr_14_eq_addr_30 and k14_needs_attention)) and (not (addr_15_eq_addr_30 and k15_needs_attention)) and (not (addr_16_eq_addr_30 and k16_needs_attention)) and (not (addr_17_eq_addr_30 and k17_needs_attention)) and (not (addr_18_eq_addr_30 and k18_needs_attention)) and (not (addr_19_eq_addr_30 and k19_needs_attention)) and (not (addr_20_eq_addr_30 and k20_needs_attention)) and (not (addr_21_eq_addr_30 and k21_needs_attention)) and (not (addr_22_eq_addr_30 and k22_needs_attention)) and (not (addr_23_eq_addr_30 and k23_needs_attention)) and (not (addr_24_eq_addr_30 and k24_needs_attention)) and (not (addr_25_eq_addr_30 and k25_needs_attention)) and (not (addr_26_eq_addr_30 and k26_needs_attention)) and (not (addr_27_eq_addr_30 and k27_needs_attention)) and (not (addr_28_eq_addr_30 and k28_needs_attention)) and (not (addr_29_eq_addr_30 and k29_needs_attention));

	k31_needs_attention <= to_bit(REQ_31) and (not (addr_0_eq_addr_31 and k0_needs_attention)) and (not (addr_1_eq_addr_31 and k1_needs_attention)) and (not (addr_2_eq_addr_31 and k2_needs_attention)) and (not (addr_3_eq_addr_31 and k3_needs_attention)) and (not (addr_4_eq_addr_31 and k4_needs_attention)) and (not (addr_5_eq_addr_31 and k5_needs_attention)) and (not (addr_6_eq_addr_31 and k6_needs_attention)) and (not (addr_7_eq_addr_31 and k7_needs_attention)) and (not (addr_8_eq_addr_31 and k8_needs_attention)) and (not (addr_9_eq_addr_31 and k9_needs_attention)) and (not (addr_10_eq_addr_31 and k10_needs_attention)) and (not (addr_11_eq_addr_31 and k11_needs_attention)) and (not (addr_12_eq_addr_31 and k12_needs_attention)) and (not (addr_13_eq_addr_31 and k13_needs_attention)) and (not (addr_14_eq_addr_31 and k14_needs_attention)) and (not (addr_15_eq_addr_31 and k15_needs_attention)) and (not (addr_16_eq_addr_31 and k16_needs_attention)) and (not (addr_17_eq_addr_31 and k17_needs_attention)) and (not (addr_18_eq_addr_31 and k18_needs_attention)) and (not (addr_19_eq_addr_31 and k19_needs_attention)) and (not (addr_20_eq_addr_31 and k20_needs_attention)) and (not (addr_21_eq_addr_31 and k21_needs_attention)) and (not (addr_22_eq_addr_31 and k22_needs_attention)) and (not (addr_23_eq_addr_31 and k23_needs_attention)) and (not (addr_24_eq_addr_31 and k24_needs_attention)) and (not (addr_25_eq_addr_31 and k25_needs_attention)) and (not (addr_26_eq_addr_31 and k26_needs_attention)) and (not (addr_27_eq_addr_31 and k27_needs_attention)) and (not (addr_28_eq_addr_31 and k28_needs_attention)) and (not (addr_29_eq_addr_31 and k29_needs_attention)) and (not (addr_30_eq_addr_31 and k30_needs_attention));


	k0_needs_bram_0 <= k0_needs_attention and not to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_1 <= k0_needs_attention and not to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_2 <= k0_needs_attention and not to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_3 <= k0_needs_attention and not to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_4 <= k0_needs_attention and not to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_5 <= k0_needs_attention and not to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_6 <= k0_needs_attention and not to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_7 <= k0_needs_attention and not to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_8 <= k0_needs_attention and     to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_9 <= k0_needs_attention and     to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_10 <= k0_needs_attention and     to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_11 <= k0_needs_attention and     to_bit(ADDR_0(12)) and not to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_12 <= k0_needs_attention and     to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_13 <= k0_needs_attention and     to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and not to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));
	k0_needs_bram_14 <= k0_needs_attention and     to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and not to_bit(ADDR_0(9));
	k0_needs_bram_15 <= k0_needs_attention and     to_bit(ADDR_0(12)) and     to_bit(ADDR_0(11)) and     to_bit(ADDR_0(10)) and     to_bit(ADDR_0(9));

	k1_needs_bram_0 <= k1_needs_attention and not to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_1 <= k1_needs_attention and not to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_2 <= k1_needs_attention and not to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_3 <= k1_needs_attention and not to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_4 <= k1_needs_attention and not to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_5 <= k1_needs_attention and not to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_6 <= k1_needs_attention and not to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_7 <= k1_needs_attention and not to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_8 <= k1_needs_attention and     to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_9 <= k1_needs_attention and     to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_10 <= k1_needs_attention and     to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_11 <= k1_needs_attention and     to_bit(ADDR_1(12)) and not to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_12 <= k1_needs_attention and     to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_13 <= k1_needs_attention and     to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and not to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));
	k1_needs_bram_14 <= k1_needs_attention and     to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and not to_bit(ADDR_1(9));
	k1_needs_bram_15 <= k1_needs_attention and     to_bit(ADDR_1(12)) and     to_bit(ADDR_1(11)) and     to_bit(ADDR_1(10)) and     to_bit(ADDR_1(9));

	k2_needs_bram_0 <= k2_needs_attention and not to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_1 <= k2_needs_attention and not to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_2 <= k2_needs_attention and not to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_3 <= k2_needs_attention and not to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_4 <= k2_needs_attention and not to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_5 <= k2_needs_attention and not to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_6 <= k2_needs_attention and not to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_7 <= k2_needs_attention and not to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_8 <= k2_needs_attention and     to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_9 <= k2_needs_attention and     to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_10 <= k2_needs_attention and     to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_11 <= k2_needs_attention and     to_bit(ADDR_2(12)) and not to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_12 <= k2_needs_attention and     to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_13 <= k2_needs_attention and     to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and not to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));
	k2_needs_bram_14 <= k2_needs_attention and     to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and not to_bit(ADDR_2(9));
	k2_needs_bram_15 <= k2_needs_attention and     to_bit(ADDR_2(12)) and     to_bit(ADDR_2(11)) and     to_bit(ADDR_2(10)) and     to_bit(ADDR_2(9));

	k3_needs_bram_0 <= k3_needs_attention and not to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_1 <= k3_needs_attention and not to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_2 <= k3_needs_attention and not to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_3 <= k3_needs_attention and not to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_4 <= k3_needs_attention and not to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_5 <= k3_needs_attention and not to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_6 <= k3_needs_attention and not to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_7 <= k3_needs_attention and not to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_8 <= k3_needs_attention and     to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_9 <= k3_needs_attention and     to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_10 <= k3_needs_attention and     to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_11 <= k3_needs_attention and     to_bit(ADDR_3(12)) and not to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_12 <= k3_needs_attention and     to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_13 <= k3_needs_attention and     to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and not to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));
	k3_needs_bram_14 <= k3_needs_attention and     to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and not to_bit(ADDR_3(9));
	k3_needs_bram_15 <= k3_needs_attention and     to_bit(ADDR_3(12)) and     to_bit(ADDR_3(11)) and     to_bit(ADDR_3(10)) and     to_bit(ADDR_3(9));

	k4_needs_bram_0 <= k4_needs_attention and not to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_1 <= k4_needs_attention and not to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_2 <= k4_needs_attention and not to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_3 <= k4_needs_attention and not to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_4 <= k4_needs_attention and not to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_5 <= k4_needs_attention and not to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_6 <= k4_needs_attention and not to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_7 <= k4_needs_attention and not to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_8 <= k4_needs_attention and     to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_9 <= k4_needs_attention and     to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_10 <= k4_needs_attention and     to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_11 <= k4_needs_attention and     to_bit(ADDR_4(12)) and not to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_12 <= k4_needs_attention and     to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_13 <= k4_needs_attention and     to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and not to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));
	k4_needs_bram_14 <= k4_needs_attention and     to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and not to_bit(ADDR_4(9));
	k4_needs_bram_15 <= k4_needs_attention and     to_bit(ADDR_4(12)) and     to_bit(ADDR_4(11)) and     to_bit(ADDR_4(10)) and     to_bit(ADDR_4(9));

	k5_needs_bram_0 <= k5_needs_attention and not to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_1 <= k5_needs_attention and not to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_2 <= k5_needs_attention and not to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_3 <= k5_needs_attention and not to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_4 <= k5_needs_attention and not to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_5 <= k5_needs_attention and not to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_6 <= k5_needs_attention and not to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_7 <= k5_needs_attention and not to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_8 <= k5_needs_attention and     to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_9 <= k5_needs_attention and     to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_10 <= k5_needs_attention and     to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_11 <= k5_needs_attention and     to_bit(ADDR_5(12)) and not to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_12 <= k5_needs_attention and     to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_13 <= k5_needs_attention and     to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and not to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));
	k5_needs_bram_14 <= k5_needs_attention and     to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and not to_bit(ADDR_5(9));
	k5_needs_bram_15 <= k5_needs_attention and     to_bit(ADDR_5(12)) and     to_bit(ADDR_5(11)) and     to_bit(ADDR_5(10)) and     to_bit(ADDR_5(9));

	k6_needs_bram_0 <= k6_needs_attention and not to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_1 <= k6_needs_attention and not to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_2 <= k6_needs_attention and not to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_3 <= k6_needs_attention and not to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_4 <= k6_needs_attention and not to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_5 <= k6_needs_attention and not to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_6 <= k6_needs_attention and not to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_7 <= k6_needs_attention and not to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_8 <= k6_needs_attention and     to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_9 <= k6_needs_attention and     to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_10 <= k6_needs_attention and     to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_11 <= k6_needs_attention and     to_bit(ADDR_6(12)) and not to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_12 <= k6_needs_attention and     to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_13 <= k6_needs_attention and     to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and not to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));
	k6_needs_bram_14 <= k6_needs_attention and     to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and not to_bit(ADDR_6(9));
	k6_needs_bram_15 <= k6_needs_attention and     to_bit(ADDR_6(12)) and     to_bit(ADDR_6(11)) and     to_bit(ADDR_6(10)) and     to_bit(ADDR_6(9));

	k7_needs_bram_0 <= k7_needs_attention and not to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_1 <= k7_needs_attention and not to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_2 <= k7_needs_attention and not to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_3 <= k7_needs_attention and not to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_4 <= k7_needs_attention and not to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_5 <= k7_needs_attention and not to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_6 <= k7_needs_attention and not to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_7 <= k7_needs_attention and not to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_8 <= k7_needs_attention and     to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_9 <= k7_needs_attention and     to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_10 <= k7_needs_attention and     to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_11 <= k7_needs_attention and     to_bit(ADDR_7(12)) and not to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_12 <= k7_needs_attention and     to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_13 <= k7_needs_attention and     to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and not to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));
	k7_needs_bram_14 <= k7_needs_attention and     to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and not to_bit(ADDR_7(9));
	k7_needs_bram_15 <= k7_needs_attention and     to_bit(ADDR_7(12)) and     to_bit(ADDR_7(11)) and     to_bit(ADDR_7(10)) and     to_bit(ADDR_7(9));

	k8_needs_bram_0 <= k8_needs_attention and not to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_1 <= k8_needs_attention and not to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_2 <= k8_needs_attention and not to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_3 <= k8_needs_attention and not to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_4 <= k8_needs_attention and not to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_5 <= k8_needs_attention and not to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_6 <= k8_needs_attention and not to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_7 <= k8_needs_attention and not to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_8 <= k8_needs_attention and     to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_9 <= k8_needs_attention and     to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_10 <= k8_needs_attention and     to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_11 <= k8_needs_attention and     to_bit(ADDR_8(12)) and not to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_12 <= k8_needs_attention and     to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_13 <= k8_needs_attention and     to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and not to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));
	k8_needs_bram_14 <= k8_needs_attention and     to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and not to_bit(ADDR_8(9));
	k8_needs_bram_15 <= k8_needs_attention and     to_bit(ADDR_8(12)) and     to_bit(ADDR_8(11)) and     to_bit(ADDR_8(10)) and     to_bit(ADDR_8(9));

	k9_needs_bram_0 <= k9_needs_attention and not to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_1 <= k9_needs_attention and not to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_2 <= k9_needs_attention and not to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_3 <= k9_needs_attention and not to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_4 <= k9_needs_attention and not to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_5 <= k9_needs_attention and not to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_6 <= k9_needs_attention and not to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_7 <= k9_needs_attention and not to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_8 <= k9_needs_attention and     to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_9 <= k9_needs_attention and     to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_10 <= k9_needs_attention and     to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_11 <= k9_needs_attention and     to_bit(ADDR_9(12)) and not to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_12 <= k9_needs_attention and     to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_13 <= k9_needs_attention and     to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and not to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));
	k9_needs_bram_14 <= k9_needs_attention and     to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and not to_bit(ADDR_9(9));
	k9_needs_bram_15 <= k9_needs_attention and     to_bit(ADDR_9(12)) and     to_bit(ADDR_9(11)) and     to_bit(ADDR_9(10)) and     to_bit(ADDR_9(9));

	k10_needs_bram_0 <= k10_needs_attention and not to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_1 <= k10_needs_attention and not to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_2 <= k10_needs_attention and not to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_3 <= k10_needs_attention and not to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_4 <= k10_needs_attention and not to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_5 <= k10_needs_attention and not to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_6 <= k10_needs_attention and not to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_7 <= k10_needs_attention and not to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_8 <= k10_needs_attention and     to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_9 <= k10_needs_attention and     to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_10 <= k10_needs_attention and     to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_11 <= k10_needs_attention and     to_bit(ADDR_10(12)) and not to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_12 <= k10_needs_attention and     to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_13 <= k10_needs_attention and     to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and not to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));
	k10_needs_bram_14 <= k10_needs_attention and     to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and not to_bit(ADDR_10(9));
	k10_needs_bram_15 <= k10_needs_attention and     to_bit(ADDR_10(12)) and     to_bit(ADDR_10(11)) and     to_bit(ADDR_10(10)) and     to_bit(ADDR_10(9));

	k11_needs_bram_0 <= k11_needs_attention and not to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_1 <= k11_needs_attention and not to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_2 <= k11_needs_attention and not to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_3 <= k11_needs_attention and not to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_4 <= k11_needs_attention and not to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_5 <= k11_needs_attention and not to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_6 <= k11_needs_attention and not to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_7 <= k11_needs_attention and not to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_8 <= k11_needs_attention and     to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_9 <= k11_needs_attention and     to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_10 <= k11_needs_attention and     to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_11 <= k11_needs_attention and     to_bit(ADDR_11(12)) and not to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_12 <= k11_needs_attention and     to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_13 <= k11_needs_attention and     to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and not to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));
	k11_needs_bram_14 <= k11_needs_attention and     to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and not to_bit(ADDR_11(9));
	k11_needs_bram_15 <= k11_needs_attention and     to_bit(ADDR_11(12)) and     to_bit(ADDR_11(11)) and     to_bit(ADDR_11(10)) and     to_bit(ADDR_11(9));

	k12_needs_bram_0 <= k12_needs_attention and not to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_1 <= k12_needs_attention and not to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_2 <= k12_needs_attention and not to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_3 <= k12_needs_attention and not to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_4 <= k12_needs_attention and not to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_5 <= k12_needs_attention and not to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_6 <= k12_needs_attention and not to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_7 <= k12_needs_attention and not to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_8 <= k12_needs_attention and     to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_9 <= k12_needs_attention and     to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_10 <= k12_needs_attention and     to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_11 <= k12_needs_attention and     to_bit(ADDR_12(12)) and not to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_12 <= k12_needs_attention and     to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_13 <= k12_needs_attention and     to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and not to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));
	k12_needs_bram_14 <= k12_needs_attention and     to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and not to_bit(ADDR_12(9));
	k12_needs_bram_15 <= k12_needs_attention and     to_bit(ADDR_12(12)) and     to_bit(ADDR_12(11)) and     to_bit(ADDR_12(10)) and     to_bit(ADDR_12(9));

	k13_needs_bram_0 <= k13_needs_attention and not to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_1 <= k13_needs_attention and not to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_2 <= k13_needs_attention and not to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_3 <= k13_needs_attention and not to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_4 <= k13_needs_attention and not to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_5 <= k13_needs_attention and not to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_6 <= k13_needs_attention and not to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_7 <= k13_needs_attention and not to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_8 <= k13_needs_attention and     to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_9 <= k13_needs_attention and     to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_10 <= k13_needs_attention and     to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_11 <= k13_needs_attention and     to_bit(ADDR_13(12)) and not to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_12 <= k13_needs_attention and     to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_13 <= k13_needs_attention and     to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and not to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));
	k13_needs_bram_14 <= k13_needs_attention and     to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and not to_bit(ADDR_13(9));
	k13_needs_bram_15 <= k13_needs_attention and     to_bit(ADDR_13(12)) and     to_bit(ADDR_13(11)) and     to_bit(ADDR_13(10)) and     to_bit(ADDR_13(9));

	k14_needs_bram_0 <= k14_needs_attention and not to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_1 <= k14_needs_attention and not to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_2 <= k14_needs_attention and not to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_3 <= k14_needs_attention and not to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_4 <= k14_needs_attention and not to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_5 <= k14_needs_attention and not to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_6 <= k14_needs_attention and not to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_7 <= k14_needs_attention and not to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_8 <= k14_needs_attention and     to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_9 <= k14_needs_attention and     to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_10 <= k14_needs_attention and     to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_11 <= k14_needs_attention and     to_bit(ADDR_14(12)) and not to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_12 <= k14_needs_attention and     to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_13 <= k14_needs_attention and     to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and not to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));
	k14_needs_bram_14 <= k14_needs_attention and     to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and not to_bit(ADDR_14(9));
	k14_needs_bram_15 <= k14_needs_attention and     to_bit(ADDR_14(12)) and     to_bit(ADDR_14(11)) and     to_bit(ADDR_14(10)) and     to_bit(ADDR_14(9));

	k15_needs_bram_0 <= k15_needs_attention and not to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_1 <= k15_needs_attention and not to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_2 <= k15_needs_attention and not to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_3 <= k15_needs_attention and not to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_4 <= k15_needs_attention and not to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_5 <= k15_needs_attention and not to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_6 <= k15_needs_attention and not to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_7 <= k15_needs_attention and not to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_8 <= k15_needs_attention and     to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_9 <= k15_needs_attention and     to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_10 <= k15_needs_attention and     to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_11 <= k15_needs_attention and     to_bit(ADDR_15(12)) and not to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_12 <= k15_needs_attention and     to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_13 <= k15_needs_attention and     to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and not to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));
	k15_needs_bram_14 <= k15_needs_attention and     to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and not to_bit(ADDR_15(9));
	k15_needs_bram_15 <= k15_needs_attention and     to_bit(ADDR_15(12)) and     to_bit(ADDR_15(11)) and     to_bit(ADDR_15(10)) and     to_bit(ADDR_15(9));

	k16_needs_bram_0 <= k16_needs_attention and not to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_1 <= k16_needs_attention and not to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_2 <= k16_needs_attention and not to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_3 <= k16_needs_attention and not to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_4 <= k16_needs_attention and not to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_5 <= k16_needs_attention and not to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_6 <= k16_needs_attention and not to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_7 <= k16_needs_attention and not to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_8 <= k16_needs_attention and     to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_9 <= k16_needs_attention and     to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_10 <= k16_needs_attention and     to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_11 <= k16_needs_attention and     to_bit(ADDR_16(12)) and not to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_12 <= k16_needs_attention and     to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_13 <= k16_needs_attention and     to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and not to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));
	k16_needs_bram_14 <= k16_needs_attention and     to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and not to_bit(ADDR_16(9));
	k16_needs_bram_15 <= k16_needs_attention and     to_bit(ADDR_16(12)) and     to_bit(ADDR_16(11)) and     to_bit(ADDR_16(10)) and     to_bit(ADDR_16(9));

	k17_needs_bram_0 <= k17_needs_attention and not to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_1 <= k17_needs_attention and not to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_2 <= k17_needs_attention and not to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_3 <= k17_needs_attention and not to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_4 <= k17_needs_attention and not to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_5 <= k17_needs_attention and not to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_6 <= k17_needs_attention and not to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_7 <= k17_needs_attention and not to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_8 <= k17_needs_attention and     to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_9 <= k17_needs_attention and     to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_10 <= k17_needs_attention and     to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_11 <= k17_needs_attention and     to_bit(ADDR_17(12)) and not to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_12 <= k17_needs_attention and     to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_13 <= k17_needs_attention and     to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and not to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));
	k17_needs_bram_14 <= k17_needs_attention and     to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and not to_bit(ADDR_17(9));
	k17_needs_bram_15 <= k17_needs_attention and     to_bit(ADDR_17(12)) and     to_bit(ADDR_17(11)) and     to_bit(ADDR_17(10)) and     to_bit(ADDR_17(9));

	k18_needs_bram_0 <= k18_needs_attention and not to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_1 <= k18_needs_attention and not to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_2 <= k18_needs_attention and not to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_3 <= k18_needs_attention and not to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_4 <= k18_needs_attention and not to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_5 <= k18_needs_attention and not to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_6 <= k18_needs_attention and not to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_7 <= k18_needs_attention and not to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_8 <= k18_needs_attention and     to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_9 <= k18_needs_attention and     to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_10 <= k18_needs_attention and     to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_11 <= k18_needs_attention and     to_bit(ADDR_18(12)) and not to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_12 <= k18_needs_attention and     to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_13 <= k18_needs_attention and     to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and not to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));
	k18_needs_bram_14 <= k18_needs_attention and     to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and not to_bit(ADDR_18(9));
	k18_needs_bram_15 <= k18_needs_attention and     to_bit(ADDR_18(12)) and     to_bit(ADDR_18(11)) and     to_bit(ADDR_18(10)) and     to_bit(ADDR_18(9));

	k19_needs_bram_0 <= k19_needs_attention and not to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_1 <= k19_needs_attention and not to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_2 <= k19_needs_attention and not to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_3 <= k19_needs_attention and not to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_4 <= k19_needs_attention and not to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_5 <= k19_needs_attention and not to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_6 <= k19_needs_attention and not to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_7 <= k19_needs_attention and not to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_8 <= k19_needs_attention and     to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_9 <= k19_needs_attention and     to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_10 <= k19_needs_attention and     to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_11 <= k19_needs_attention and     to_bit(ADDR_19(12)) and not to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_12 <= k19_needs_attention and     to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_13 <= k19_needs_attention and     to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and not to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));
	k19_needs_bram_14 <= k19_needs_attention and     to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and not to_bit(ADDR_19(9));
	k19_needs_bram_15 <= k19_needs_attention and     to_bit(ADDR_19(12)) and     to_bit(ADDR_19(11)) and     to_bit(ADDR_19(10)) and     to_bit(ADDR_19(9));

	k20_needs_bram_0 <= k20_needs_attention and not to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_1 <= k20_needs_attention and not to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_2 <= k20_needs_attention and not to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_3 <= k20_needs_attention and not to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_4 <= k20_needs_attention and not to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_5 <= k20_needs_attention and not to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_6 <= k20_needs_attention and not to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_7 <= k20_needs_attention and not to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_8 <= k20_needs_attention and     to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_9 <= k20_needs_attention and     to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_10 <= k20_needs_attention and     to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_11 <= k20_needs_attention and     to_bit(ADDR_20(12)) and not to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_12 <= k20_needs_attention and     to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_13 <= k20_needs_attention and     to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and not to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));
	k20_needs_bram_14 <= k20_needs_attention and     to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and not to_bit(ADDR_20(9));
	k20_needs_bram_15 <= k20_needs_attention and     to_bit(ADDR_20(12)) and     to_bit(ADDR_20(11)) and     to_bit(ADDR_20(10)) and     to_bit(ADDR_20(9));

	k21_needs_bram_0 <= k21_needs_attention and not to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_1 <= k21_needs_attention and not to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_2 <= k21_needs_attention and not to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_3 <= k21_needs_attention and not to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_4 <= k21_needs_attention and not to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_5 <= k21_needs_attention and not to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_6 <= k21_needs_attention and not to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_7 <= k21_needs_attention and not to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_8 <= k21_needs_attention and     to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_9 <= k21_needs_attention and     to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_10 <= k21_needs_attention and     to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_11 <= k21_needs_attention and     to_bit(ADDR_21(12)) and not to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_12 <= k21_needs_attention and     to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_13 <= k21_needs_attention and     to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and not to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));
	k21_needs_bram_14 <= k21_needs_attention and     to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and not to_bit(ADDR_21(9));
	k21_needs_bram_15 <= k21_needs_attention and     to_bit(ADDR_21(12)) and     to_bit(ADDR_21(11)) and     to_bit(ADDR_21(10)) and     to_bit(ADDR_21(9));

	k22_needs_bram_0 <= k22_needs_attention and not to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_1 <= k22_needs_attention and not to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_2 <= k22_needs_attention and not to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_3 <= k22_needs_attention and not to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_4 <= k22_needs_attention and not to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_5 <= k22_needs_attention and not to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_6 <= k22_needs_attention and not to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_7 <= k22_needs_attention and not to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_8 <= k22_needs_attention and     to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_9 <= k22_needs_attention and     to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_10 <= k22_needs_attention and     to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_11 <= k22_needs_attention and     to_bit(ADDR_22(12)) and not to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_12 <= k22_needs_attention and     to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_13 <= k22_needs_attention and     to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and not to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));
	k22_needs_bram_14 <= k22_needs_attention and     to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and not to_bit(ADDR_22(9));
	k22_needs_bram_15 <= k22_needs_attention and     to_bit(ADDR_22(12)) and     to_bit(ADDR_22(11)) and     to_bit(ADDR_22(10)) and     to_bit(ADDR_22(9));

	k23_needs_bram_0 <= k23_needs_attention and not to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_1 <= k23_needs_attention and not to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_2 <= k23_needs_attention and not to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_3 <= k23_needs_attention and not to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_4 <= k23_needs_attention and not to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_5 <= k23_needs_attention and not to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_6 <= k23_needs_attention and not to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_7 <= k23_needs_attention and not to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_8 <= k23_needs_attention and     to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_9 <= k23_needs_attention and     to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_10 <= k23_needs_attention and     to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_11 <= k23_needs_attention and     to_bit(ADDR_23(12)) and not to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_12 <= k23_needs_attention and     to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_13 <= k23_needs_attention and     to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and not to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));
	k23_needs_bram_14 <= k23_needs_attention and     to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and not to_bit(ADDR_23(9));
	k23_needs_bram_15 <= k23_needs_attention and     to_bit(ADDR_23(12)) and     to_bit(ADDR_23(11)) and     to_bit(ADDR_23(10)) and     to_bit(ADDR_23(9));

	k24_needs_bram_0 <= k24_needs_attention and not to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_1 <= k24_needs_attention and not to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_2 <= k24_needs_attention and not to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_3 <= k24_needs_attention and not to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_4 <= k24_needs_attention and not to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_5 <= k24_needs_attention and not to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_6 <= k24_needs_attention and not to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_7 <= k24_needs_attention and not to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_8 <= k24_needs_attention and     to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_9 <= k24_needs_attention and     to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_10 <= k24_needs_attention and     to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_11 <= k24_needs_attention and     to_bit(ADDR_24(12)) and not to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_12 <= k24_needs_attention and     to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_13 <= k24_needs_attention and     to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and not to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));
	k24_needs_bram_14 <= k24_needs_attention and     to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and not to_bit(ADDR_24(9));
	k24_needs_bram_15 <= k24_needs_attention and     to_bit(ADDR_24(12)) and     to_bit(ADDR_24(11)) and     to_bit(ADDR_24(10)) and     to_bit(ADDR_24(9));

	k25_needs_bram_0 <= k25_needs_attention and not to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_1 <= k25_needs_attention and not to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_2 <= k25_needs_attention and not to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_3 <= k25_needs_attention and not to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_4 <= k25_needs_attention and not to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_5 <= k25_needs_attention and not to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_6 <= k25_needs_attention and not to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_7 <= k25_needs_attention and not to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_8 <= k25_needs_attention and     to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_9 <= k25_needs_attention and     to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_10 <= k25_needs_attention and     to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_11 <= k25_needs_attention and     to_bit(ADDR_25(12)) and not to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_12 <= k25_needs_attention and     to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_13 <= k25_needs_attention and     to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and not to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));
	k25_needs_bram_14 <= k25_needs_attention and     to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and not to_bit(ADDR_25(9));
	k25_needs_bram_15 <= k25_needs_attention and     to_bit(ADDR_25(12)) and     to_bit(ADDR_25(11)) and     to_bit(ADDR_25(10)) and     to_bit(ADDR_25(9));

	k26_needs_bram_0 <= k26_needs_attention and not to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_1 <= k26_needs_attention and not to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_2 <= k26_needs_attention and not to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_3 <= k26_needs_attention and not to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_4 <= k26_needs_attention and not to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_5 <= k26_needs_attention and not to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_6 <= k26_needs_attention and not to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_7 <= k26_needs_attention and not to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_8 <= k26_needs_attention and     to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_9 <= k26_needs_attention and     to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_10 <= k26_needs_attention and     to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_11 <= k26_needs_attention and     to_bit(ADDR_26(12)) and not to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_12 <= k26_needs_attention and     to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_13 <= k26_needs_attention and     to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and not to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));
	k26_needs_bram_14 <= k26_needs_attention and     to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and not to_bit(ADDR_26(9));
	k26_needs_bram_15 <= k26_needs_attention and     to_bit(ADDR_26(12)) and     to_bit(ADDR_26(11)) and     to_bit(ADDR_26(10)) and     to_bit(ADDR_26(9));

	k27_needs_bram_0 <= k27_needs_attention and not to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_1 <= k27_needs_attention and not to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_2 <= k27_needs_attention and not to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_3 <= k27_needs_attention and not to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_4 <= k27_needs_attention and not to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_5 <= k27_needs_attention and not to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_6 <= k27_needs_attention and not to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_7 <= k27_needs_attention and not to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_8 <= k27_needs_attention and     to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_9 <= k27_needs_attention and     to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_10 <= k27_needs_attention and     to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_11 <= k27_needs_attention and     to_bit(ADDR_27(12)) and not to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_12 <= k27_needs_attention and     to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_13 <= k27_needs_attention and     to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and not to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));
	k27_needs_bram_14 <= k27_needs_attention and     to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and not to_bit(ADDR_27(9));
	k27_needs_bram_15 <= k27_needs_attention and     to_bit(ADDR_27(12)) and     to_bit(ADDR_27(11)) and     to_bit(ADDR_27(10)) and     to_bit(ADDR_27(9));

	k28_needs_bram_0 <= k28_needs_attention and not to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_1 <= k28_needs_attention and not to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_2 <= k28_needs_attention and not to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_3 <= k28_needs_attention and not to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_4 <= k28_needs_attention and not to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_5 <= k28_needs_attention and not to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_6 <= k28_needs_attention and not to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_7 <= k28_needs_attention and not to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_8 <= k28_needs_attention and     to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_9 <= k28_needs_attention and     to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_10 <= k28_needs_attention and     to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_11 <= k28_needs_attention and     to_bit(ADDR_28(12)) and not to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_12 <= k28_needs_attention and     to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_13 <= k28_needs_attention and     to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and not to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));
	k28_needs_bram_14 <= k28_needs_attention and     to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and not to_bit(ADDR_28(9));
	k28_needs_bram_15 <= k28_needs_attention and     to_bit(ADDR_28(12)) and     to_bit(ADDR_28(11)) and     to_bit(ADDR_28(10)) and     to_bit(ADDR_28(9));

	k29_needs_bram_0 <= k29_needs_attention and not to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_1 <= k29_needs_attention and not to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_2 <= k29_needs_attention and not to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_3 <= k29_needs_attention and not to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_4 <= k29_needs_attention and not to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_5 <= k29_needs_attention and not to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_6 <= k29_needs_attention and not to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_7 <= k29_needs_attention and not to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_8 <= k29_needs_attention and     to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_9 <= k29_needs_attention and     to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_10 <= k29_needs_attention and     to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_11 <= k29_needs_attention and     to_bit(ADDR_29(12)) and not to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_12 <= k29_needs_attention and     to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_13 <= k29_needs_attention and     to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and not to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));
	k29_needs_bram_14 <= k29_needs_attention and     to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and not to_bit(ADDR_29(9));
	k29_needs_bram_15 <= k29_needs_attention and     to_bit(ADDR_29(12)) and     to_bit(ADDR_29(11)) and     to_bit(ADDR_29(10)) and     to_bit(ADDR_29(9));

	k30_needs_bram_0 <= k30_needs_attention and not to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_1 <= k30_needs_attention and not to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_2 <= k30_needs_attention and not to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_3 <= k30_needs_attention and not to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_4 <= k30_needs_attention and not to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_5 <= k30_needs_attention and not to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_6 <= k30_needs_attention and not to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_7 <= k30_needs_attention and not to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_8 <= k30_needs_attention and     to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_9 <= k30_needs_attention and     to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_10 <= k30_needs_attention and     to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_11 <= k30_needs_attention and     to_bit(ADDR_30(12)) and not to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_12 <= k30_needs_attention and     to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_13 <= k30_needs_attention and     to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and not to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));
	k30_needs_bram_14 <= k30_needs_attention and     to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and not to_bit(ADDR_30(9));
	k30_needs_bram_15 <= k30_needs_attention and     to_bit(ADDR_30(12)) and     to_bit(ADDR_30(11)) and     to_bit(ADDR_30(10)) and     to_bit(ADDR_30(9));

	k31_needs_bram_0 <= k31_needs_attention and not to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_1 <= k31_needs_attention and not to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_2 <= k31_needs_attention and not to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_3 <= k31_needs_attention and not to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_4 <= k31_needs_attention and not to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_5 <= k31_needs_attention and not to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_6 <= k31_needs_attention and not to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_7 <= k31_needs_attention and not to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_8 <= k31_needs_attention and     to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_9 <= k31_needs_attention and     to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_10 <= k31_needs_attention and     to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_11 <= k31_needs_attention and     to_bit(ADDR_31(12)) and not to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_12 <= k31_needs_attention and     to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_13 <= k31_needs_attention and     to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and not to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));
	k31_needs_bram_14 <= k31_needs_attention and     to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and not to_bit(ADDR_31(9));
	k31_needs_bram_15 <= k31_needs_attention and     to_bit(ADDR_31(12)) and     to_bit(ADDR_31(11)) and     to_bit(ADDR_31(10)) and     to_bit(ADDR_31(9));


	bram_0_input_sel(4) <= not ((k0_needs_bram_0 or k1_needs_bram_0 or k2_needs_bram_0 or k3_needs_bram_0 or k4_needs_bram_0 or k5_needs_bram_0 or k6_needs_bram_0 or k7_needs_bram_0 or k8_needs_bram_0 or k9_needs_bram_0 or k10_needs_bram_0 or k11_needs_bram_0 or k12_needs_bram_0 or k13_needs_bram_0 or k14_needs_bram_0 or k15_needs_bram_0));
	bram_2_input_sel(4) <= not ((k0_needs_bram_1 or k1_needs_bram_1 or k2_needs_bram_1 or k3_needs_bram_1 or k4_needs_bram_1 or k5_needs_bram_1 or k6_needs_bram_1 or k7_needs_bram_1 or k8_needs_bram_1 or k9_needs_bram_1 or k10_needs_bram_1 or k11_needs_bram_1 or k12_needs_bram_1 or k13_needs_bram_1 or k14_needs_bram_1 or k15_needs_bram_1));
	bram_4_input_sel(4) <= not ((k0_needs_bram_2 or k1_needs_bram_2 or k2_needs_bram_2 or k3_needs_bram_2 or k4_needs_bram_2 or k5_needs_bram_2 or k6_needs_bram_2 or k7_needs_bram_2 or k8_needs_bram_2 or k9_needs_bram_2 or k10_needs_bram_2 or k11_needs_bram_2 or k12_needs_bram_2 or k13_needs_bram_2 or k14_needs_bram_2 or k15_needs_bram_2));
	bram_6_input_sel(4) <= not ((k0_needs_bram_3 or k1_needs_bram_3 or k2_needs_bram_3 or k3_needs_bram_3 or k4_needs_bram_3 or k5_needs_bram_3 or k6_needs_bram_3 or k7_needs_bram_3 or k8_needs_bram_3 or k9_needs_bram_3 or k10_needs_bram_3 or k11_needs_bram_3 or k12_needs_bram_3 or k13_needs_bram_3 or k14_needs_bram_3 or k15_needs_bram_3));
	bram_8_input_sel(4) <= not ((k0_needs_bram_4 or k1_needs_bram_4 or k2_needs_bram_4 or k3_needs_bram_4 or k4_needs_bram_4 or k5_needs_bram_4 or k6_needs_bram_4 or k7_needs_bram_4 or k8_needs_bram_4 or k9_needs_bram_4 or k10_needs_bram_4 or k11_needs_bram_4 or k12_needs_bram_4 or k13_needs_bram_4 or k14_needs_bram_4 or k15_needs_bram_4));
	bram_10_input_sel(4) <= not ((k0_needs_bram_5 or k1_needs_bram_5 or k2_needs_bram_5 or k3_needs_bram_5 or k4_needs_bram_5 or k5_needs_bram_5 or k6_needs_bram_5 or k7_needs_bram_5 or k8_needs_bram_5 or k9_needs_bram_5 or k10_needs_bram_5 or k11_needs_bram_5 or k12_needs_bram_5 or k13_needs_bram_5 or k14_needs_bram_5 or k15_needs_bram_5));
	bram_12_input_sel(4) <= not ((k0_needs_bram_6 or k1_needs_bram_6 or k2_needs_bram_6 or k3_needs_bram_6 or k4_needs_bram_6 or k5_needs_bram_6 or k6_needs_bram_6 or k7_needs_bram_6 or k8_needs_bram_6 or k9_needs_bram_6 or k10_needs_bram_6 or k11_needs_bram_6 or k12_needs_bram_6 or k13_needs_bram_6 or k14_needs_bram_6 or k15_needs_bram_6));
	bram_14_input_sel(4) <= not ((k0_needs_bram_7 or k1_needs_bram_7 or k2_needs_bram_7 or k3_needs_bram_7 or k4_needs_bram_7 or k5_needs_bram_7 or k6_needs_bram_7 or k7_needs_bram_7 or k8_needs_bram_7 or k9_needs_bram_7 or k10_needs_bram_7 or k11_needs_bram_7 or k12_needs_bram_7 or k13_needs_bram_7 or k14_needs_bram_7 or k15_needs_bram_7));
	bram_16_input_sel(4) <= not ((k0_needs_bram_8 or k1_needs_bram_8 or k2_needs_bram_8 or k3_needs_bram_8 or k4_needs_bram_8 or k5_needs_bram_8 or k6_needs_bram_8 or k7_needs_bram_8 or k8_needs_bram_8 or k9_needs_bram_8 or k10_needs_bram_8 or k11_needs_bram_8 or k12_needs_bram_8 or k13_needs_bram_8 or k14_needs_bram_8 or k15_needs_bram_8));
	bram_18_input_sel(4) <= not ((k0_needs_bram_9 or k1_needs_bram_9 or k2_needs_bram_9 or k3_needs_bram_9 or k4_needs_bram_9 or k5_needs_bram_9 or k6_needs_bram_9 or k7_needs_bram_9 or k8_needs_bram_9 or k9_needs_bram_9 or k10_needs_bram_9 or k11_needs_bram_9 or k12_needs_bram_9 or k13_needs_bram_9 or k14_needs_bram_9 or k15_needs_bram_9));
	bram_20_input_sel(4) <= not ((k0_needs_bram_10 or k1_needs_bram_10 or k2_needs_bram_10 or k3_needs_bram_10 or k4_needs_bram_10 or k5_needs_bram_10 or k6_needs_bram_10 or k7_needs_bram_10 or k8_needs_bram_10 or k9_needs_bram_10 or k10_needs_bram_10 or k11_needs_bram_10 or k12_needs_bram_10 or k13_needs_bram_10 or k14_needs_bram_10 or k15_needs_bram_10));
	bram_22_input_sel(4) <= not ((k0_needs_bram_11 or k1_needs_bram_11 or k2_needs_bram_11 or k3_needs_bram_11 or k4_needs_bram_11 or k5_needs_bram_11 or k6_needs_bram_11 or k7_needs_bram_11 or k8_needs_bram_11 or k9_needs_bram_11 or k10_needs_bram_11 or k11_needs_bram_11 or k12_needs_bram_11 or k13_needs_bram_11 or k14_needs_bram_11 or k15_needs_bram_11));
	bram_24_input_sel(4) <= not ((k0_needs_bram_12 or k1_needs_bram_12 or k2_needs_bram_12 or k3_needs_bram_12 or k4_needs_bram_12 or k5_needs_bram_12 or k6_needs_bram_12 or k7_needs_bram_12 or k8_needs_bram_12 or k9_needs_bram_12 or k10_needs_bram_12 or k11_needs_bram_12 or k12_needs_bram_12 or k13_needs_bram_12 or k14_needs_bram_12 or k15_needs_bram_12));
	bram_26_input_sel(4) <= not ((k0_needs_bram_13 or k1_needs_bram_13 or k2_needs_bram_13 or k3_needs_bram_13 or k4_needs_bram_13 or k5_needs_bram_13 or k6_needs_bram_13 or k7_needs_bram_13 or k8_needs_bram_13 or k9_needs_bram_13 or k10_needs_bram_13 or k11_needs_bram_13 or k12_needs_bram_13 or k13_needs_bram_13 or k14_needs_bram_13 or k15_needs_bram_13));
	bram_28_input_sel(4) <= not ((k0_needs_bram_14 or k1_needs_bram_14 or k2_needs_bram_14 or k3_needs_bram_14 or k4_needs_bram_14 or k5_needs_bram_14 or k6_needs_bram_14 or k7_needs_bram_14 or k8_needs_bram_14 or k9_needs_bram_14 or k10_needs_bram_14 or k11_needs_bram_14 or k12_needs_bram_14 or k13_needs_bram_14 or k14_needs_bram_14 or k15_needs_bram_14));
	bram_30_input_sel(4) <= not ((k0_needs_bram_15 or k1_needs_bram_15 or k2_needs_bram_15 or k3_needs_bram_15 or k4_needs_bram_15 or k5_needs_bram_15 or k6_needs_bram_15 or k7_needs_bram_15 or k8_needs_bram_15 or k9_needs_bram_15 or k10_needs_bram_15 or k11_needs_bram_15 or k12_needs_bram_15 or k13_needs_bram_15 or k14_needs_bram_15 or k15_needs_bram_15));

	bram_0_input_sel(3) <= not ((k0_needs_bram_0 or k1_needs_bram_0 or k2_needs_bram_0 or k3_needs_bram_0 or k4_needs_bram_0 or k5_needs_bram_0 or k6_needs_bram_0 or k7_needs_bram_0) or ((k16_needs_bram_0 or k17_needs_bram_0 or k18_needs_bram_0 or k19_needs_bram_0 or k20_needs_bram_0 or k21_needs_bram_0 or k22_needs_bram_0 or k23_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0) and (not k13_needs_bram_0) and (not k12_needs_bram_0) and (not k11_needs_bram_0) and (not k10_needs_bram_0) and (not k9_needs_bram_0) and (not k8_needs_bram_0)));
	bram_2_input_sel(3) <= not ((k0_needs_bram_1 or k1_needs_bram_1 or k2_needs_bram_1 or k3_needs_bram_1 or k4_needs_bram_1 or k5_needs_bram_1 or k6_needs_bram_1 or k7_needs_bram_1) or ((k16_needs_bram_1 or k17_needs_bram_1 or k18_needs_bram_1 or k19_needs_bram_1 or k20_needs_bram_1 or k21_needs_bram_1 or k22_needs_bram_1 or k23_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1) and (not k13_needs_bram_1) and (not k12_needs_bram_1) and (not k11_needs_bram_1) and (not k10_needs_bram_1) and (not k9_needs_bram_1) and (not k8_needs_bram_1)));
	bram_4_input_sel(3) <= not ((k0_needs_bram_2 or k1_needs_bram_2 or k2_needs_bram_2 or k3_needs_bram_2 or k4_needs_bram_2 or k5_needs_bram_2 or k6_needs_bram_2 or k7_needs_bram_2) or ((k16_needs_bram_2 or k17_needs_bram_2 or k18_needs_bram_2 or k19_needs_bram_2 or k20_needs_bram_2 or k21_needs_bram_2 or k22_needs_bram_2 or k23_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2) and (not k13_needs_bram_2) and (not k12_needs_bram_2) and (not k11_needs_bram_2) and (not k10_needs_bram_2) and (not k9_needs_bram_2) and (not k8_needs_bram_2)));
	bram_6_input_sel(3) <= not ((k0_needs_bram_3 or k1_needs_bram_3 or k2_needs_bram_3 or k3_needs_bram_3 or k4_needs_bram_3 or k5_needs_bram_3 or k6_needs_bram_3 or k7_needs_bram_3) or ((k16_needs_bram_3 or k17_needs_bram_3 or k18_needs_bram_3 or k19_needs_bram_3 or k20_needs_bram_3 or k21_needs_bram_3 or k22_needs_bram_3 or k23_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3) and (not k13_needs_bram_3) and (not k12_needs_bram_3) and (not k11_needs_bram_3) and (not k10_needs_bram_3) and (not k9_needs_bram_3) and (not k8_needs_bram_3)));
	bram_8_input_sel(3) <= not ((k0_needs_bram_4 or k1_needs_bram_4 or k2_needs_bram_4 or k3_needs_bram_4 or k4_needs_bram_4 or k5_needs_bram_4 or k6_needs_bram_4 or k7_needs_bram_4) or ((k16_needs_bram_4 or k17_needs_bram_4 or k18_needs_bram_4 or k19_needs_bram_4 or k20_needs_bram_4 or k21_needs_bram_4 or k22_needs_bram_4 or k23_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4) and (not k13_needs_bram_4) and (not k12_needs_bram_4) and (not k11_needs_bram_4) and (not k10_needs_bram_4) and (not k9_needs_bram_4) and (not k8_needs_bram_4)));
	bram_10_input_sel(3) <= not ((k0_needs_bram_5 or k1_needs_bram_5 or k2_needs_bram_5 or k3_needs_bram_5 or k4_needs_bram_5 or k5_needs_bram_5 or k6_needs_bram_5 or k7_needs_bram_5) or ((k16_needs_bram_5 or k17_needs_bram_5 or k18_needs_bram_5 or k19_needs_bram_5 or k20_needs_bram_5 or k21_needs_bram_5 or k22_needs_bram_5 or k23_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5) and (not k13_needs_bram_5) and (not k12_needs_bram_5) and (not k11_needs_bram_5) and (not k10_needs_bram_5) and (not k9_needs_bram_5) and (not k8_needs_bram_5)));
	bram_12_input_sel(3) <= not ((k0_needs_bram_6 or k1_needs_bram_6 or k2_needs_bram_6 or k3_needs_bram_6 or k4_needs_bram_6 or k5_needs_bram_6 or k6_needs_bram_6 or k7_needs_bram_6) or ((k16_needs_bram_6 or k17_needs_bram_6 or k18_needs_bram_6 or k19_needs_bram_6 or k20_needs_bram_6 or k21_needs_bram_6 or k22_needs_bram_6 or k23_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6) and (not k13_needs_bram_6) and (not k12_needs_bram_6) and (not k11_needs_bram_6) and (not k10_needs_bram_6) and (not k9_needs_bram_6) and (not k8_needs_bram_6)));
	bram_14_input_sel(3) <= not ((k0_needs_bram_7 or k1_needs_bram_7 or k2_needs_bram_7 or k3_needs_bram_7 or k4_needs_bram_7 or k5_needs_bram_7 or k6_needs_bram_7 or k7_needs_bram_7) or ((k16_needs_bram_7 or k17_needs_bram_7 or k18_needs_bram_7 or k19_needs_bram_7 or k20_needs_bram_7 or k21_needs_bram_7 or k22_needs_bram_7 or k23_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7) and (not k13_needs_bram_7) and (not k12_needs_bram_7) and (not k11_needs_bram_7) and (not k10_needs_bram_7) and (not k9_needs_bram_7) and (not k8_needs_bram_7)));
	bram_16_input_sel(3) <= not ((k0_needs_bram_8 or k1_needs_bram_8 or k2_needs_bram_8 or k3_needs_bram_8 or k4_needs_bram_8 or k5_needs_bram_8 or k6_needs_bram_8 or k7_needs_bram_8) or ((k16_needs_bram_8 or k17_needs_bram_8 or k18_needs_bram_8 or k19_needs_bram_8 or k20_needs_bram_8 or k21_needs_bram_8 or k22_needs_bram_8 or k23_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8) and (not k13_needs_bram_8) and (not k12_needs_bram_8) and (not k11_needs_bram_8) and (not k10_needs_bram_8) and (not k9_needs_bram_8) and (not k8_needs_bram_8)));
	bram_18_input_sel(3) <= not ((k0_needs_bram_9 or k1_needs_bram_9 or k2_needs_bram_9 or k3_needs_bram_9 or k4_needs_bram_9 or k5_needs_bram_9 or k6_needs_bram_9 or k7_needs_bram_9) or ((k16_needs_bram_9 or k17_needs_bram_9 or k18_needs_bram_9 or k19_needs_bram_9 or k20_needs_bram_9 or k21_needs_bram_9 or k22_needs_bram_9 or k23_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9) and (not k13_needs_bram_9) and (not k12_needs_bram_9) and (not k11_needs_bram_9) and (not k10_needs_bram_9) and (not k9_needs_bram_9) and (not k8_needs_bram_9)));
	bram_20_input_sel(3) <= not ((k0_needs_bram_10 or k1_needs_bram_10 or k2_needs_bram_10 or k3_needs_bram_10 or k4_needs_bram_10 or k5_needs_bram_10 or k6_needs_bram_10 or k7_needs_bram_10) or ((k16_needs_bram_10 or k17_needs_bram_10 or k18_needs_bram_10 or k19_needs_bram_10 or k20_needs_bram_10 or k21_needs_bram_10 or k22_needs_bram_10 or k23_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10) and (not k13_needs_bram_10) and (not k12_needs_bram_10) and (not k11_needs_bram_10) and (not k10_needs_bram_10) and (not k9_needs_bram_10) and (not k8_needs_bram_10)));
	bram_22_input_sel(3) <= not ((k0_needs_bram_11 or k1_needs_bram_11 or k2_needs_bram_11 or k3_needs_bram_11 or k4_needs_bram_11 or k5_needs_bram_11 or k6_needs_bram_11 or k7_needs_bram_11) or ((k16_needs_bram_11 or k17_needs_bram_11 or k18_needs_bram_11 or k19_needs_bram_11 or k20_needs_bram_11 or k21_needs_bram_11 or k22_needs_bram_11 or k23_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11) and (not k13_needs_bram_11) and (not k12_needs_bram_11) and (not k11_needs_bram_11) and (not k10_needs_bram_11) and (not k9_needs_bram_11) and (not k8_needs_bram_11)));
	bram_24_input_sel(3) <= not ((k0_needs_bram_12 or k1_needs_bram_12 or k2_needs_bram_12 or k3_needs_bram_12 or k4_needs_bram_12 or k5_needs_bram_12 or k6_needs_bram_12 or k7_needs_bram_12) or ((k16_needs_bram_12 or k17_needs_bram_12 or k18_needs_bram_12 or k19_needs_bram_12 or k20_needs_bram_12 or k21_needs_bram_12 or k22_needs_bram_12 or k23_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12) and (not k13_needs_bram_12) and (not k12_needs_bram_12) and (not k11_needs_bram_12) and (not k10_needs_bram_12) and (not k9_needs_bram_12) and (not k8_needs_bram_12)));
	bram_26_input_sel(3) <= not ((k0_needs_bram_13 or k1_needs_bram_13 or k2_needs_bram_13 or k3_needs_bram_13 or k4_needs_bram_13 or k5_needs_bram_13 or k6_needs_bram_13 or k7_needs_bram_13) or ((k16_needs_bram_13 or k17_needs_bram_13 or k18_needs_bram_13 or k19_needs_bram_13 or k20_needs_bram_13 or k21_needs_bram_13 or k22_needs_bram_13 or k23_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13) and (not k13_needs_bram_13) and (not k12_needs_bram_13) and (not k11_needs_bram_13) and (not k10_needs_bram_13) and (not k9_needs_bram_13) and (not k8_needs_bram_13)));
	bram_28_input_sel(3) <= not ((k0_needs_bram_14 or k1_needs_bram_14 or k2_needs_bram_14 or k3_needs_bram_14 or k4_needs_bram_14 or k5_needs_bram_14 or k6_needs_bram_14 or k7_needs_bram_14) or ((k16_needs_bram_14 or k17_needs_bram_14 or k18_needs_bram_14 or k19_needs_bram_14 or k20_needs_bram_14 or k21_needs_bram_14 or k22_needs_bram_14 or k23_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14) and (not k13_needs_bram_14) and (not k12_needs_bram_14) and (not k11_needs_bram_14) and (not k10_needs_bram_14) and (not k9_needs_bram_14) and (not k8_needs_bram_14)));
	bram_30_input_sel(3) <= not ((k0_needs_bram_15 or k1_needs_bram_15 or k2_needs_bram_15 or k3_needs_bram_15 or k4_needs_bram_15 or k5_needs_bram_15 or k6_needs_bram_15 or k7_needs_bram_15) or ((k16_needs_bram_15 or k17_needs_bram_15 or k18_needs_bram_15 or k19_needs_bram_15 or k20_needs_bram_15 or k21_needs_bram_15 or k22_needs_bram_15 or k23_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15) and (not k13_needs_bram_15) and (not k12_needs_bram_15) and (not k11_needs_bram_15) and (not k10_needs_bram_15) and (not k9_needs_bram_15) and (not k8_needs_bram_15)));

	bram_0_input_sel(2) <= not ((k0_needs_bram_0 or k1_needs_bram_0 or k2_needs_bram_0 or k3_needs_bram_0) or ((k8_needs_bram_0 or k9_needs_bram_0 or k10_needs_bram_0 or k11_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k5_needs_bram_0) and (not k4_needs_bram_0)) or ((k16_needs_bram_0 or k17_needs_bram_0 or k18_needs_bram_0 or k19_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k5_needs_bram_0) and (not k4_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0) and (not k13_needs_bram_0) and (not k12_needs_bram_0)) or ((k24_needs_bram_0 or k25_needs_bram_0 or k26_needs_bram_0 or k27_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k5_needs_bram_0) and (not k4_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0) and (not k13_needs_bram_0) and (not k12_needs_bram_0) and (not k23_needs_bram_0) and (not k22_needs_bram_0) and (not k21_needs_bram_0) and (not k20_needs_bram_0)));
	bram_2_input_sel(2) <= not ((k0_needs_bram_1 or k1_needs_bram_1 or k2_needs_bram_1 or k3_needs_bram_1) or ((k8_needs_bram_1 or k9_needs_bram_1 or k10_needs_bram_1 or k11_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k5_needs_bram_1) and (not k4_needs_bram_1)) or ((k16_needs_bram_1 or k17_needs_bram_1 or k18_needs_bram_1 or k19_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k5_needs_bram_1) and (not k4_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1) and (not k13_needs_bram_1) and (not k12_needs_bram_1)) or ((k24_needs_bram_1 or k25_needs_bram_1 or k26_needs_bram_1 or k27_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k5_needs_bram_1) and (not k4_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1) and (not k13_needs_bram_1) and (not k12_needs_bram_1) and (not k23_needs_bram_1) and (not k22_needs_bram_1) and (not k21_needs_bram_1) and (not k20_needs_bram_1)));
	bram_4_input_sel(2) <= not ((k0_needs_bram_2 or k1_needs_bram_2 or k2_needs_bram_2 or k3_needs_bram_2) or ((k8_needs_bram_2 or k9_needs_bram_2 or k10_needs_bram_2 or k11_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k5_needs_bram_2) and (not k4_needs_bram_2)) or ((k16_needs_bram_2 or k17_needs_bram_2 or k18_needs_bram_2 or k19_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k5_needs_bram_2) and (not k4_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2) and (not k13_needs_bram_2) and (not k12_needs_bram_2)) or ((k24_needs_bram_2 or k25_needs_bram_2 or k26_needs_bram_2 or k27_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k5_needs_bram_2) and (not k4_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2) and (not k13_needs_bram_2) and (not k12_needs_bram_2) and (not k23_needs_bram_2) and (not k22_needs_bram_2) and (not k21_needs_bram_2) and (not k20_needs_bram_2)));
	bram_6_input_sel(2) <= not ((k0_needs_bram_3 or k1_needs_bram_3 or k2_needs_bram_3 or k3_needs_bram_3) or ((k8_needs_bram_3 or k9_needs_bram_3 or k10_needs_bram_3 or k11_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k5_needs_bram_3) and (not k4_needs_bram_3)) or ((k16_needs_bram_3 or k17_needs_bram_3 or k18_needs_bram_3 or k19_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k5_needs_bram_3) and (not k4_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3) and (not k13_needs_bram_3) and (not k12_needs_bram_3)) or ((k24_needs_bram_3 or k25_needs_bram_3 or k26_needs_bram_3 or k27_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k5_needs_bram_3) and (not k4_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3) and (not k13_needs_bram_3) and (not k12_needs_bram_3) and (not k23_needs_bram_3) and (not k22_needs_bram_3) and (not k21_needs_bram_3) and (not k20_needs_bram_3)));
	bram_8_input_sel(2) <= not ((k0_needs_bram_4 or k1_needs_bram_4 or k2_needs_bram_4 or k3_needs_bram_4) or ((k8_needs_bram_4 or k9_needs_bram_4 or k10_needs_bram_4 or k11_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k5_needs_bram_4) and (not k4_needs_bram_4)) or ((k16_needs_bram_4 or k17_needs_bram_4 or k18_needs_bram_4 or k19_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k5_needs_bram_4) and (not k4_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4) and (not k13_needs_bram_4) and (not k12_needs_bram_4)) or ((k24_needs_bram_4 or k25_needs_bram_4 or k26_needs_bram_4 or k27_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k5_needs_bram_4) and (not k4_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4) and (not k13_needs_bram_4) and (not k12_needs_bram_4) and (not k23_needs_bram_4) and (not k22_needs_bram_4) and (not k21_needs_bram_4) and (not k20_needs_bram_4)));
	bram_10_input_sel(2) <= not ((k0_needs_bram_5 or k1_needs_bram_5 or k2_needs_bram_5 or k3_needs_bram_5) or ((k8_needs_bram_5 or k9_needs_bram_5 or k10_needs_bram_5 or k11_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k5_needs_bram_5) and (not k4_needs_bram_5)) or ((k16_needs_bram_5 or k17_needs_bram_5 or k18_needs_bram_5 or k19_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k5_needs_bram_5) and (not k4_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5) and (not k13_needs_bram_5) and (not k12_needs_bram_5)) or ((k24_needs_bram_5 or k25_needs_bram_5 or k26_needs_bram_5 or k27_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k5_needs_bram_5) and (not k4_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5) and (not k13_needs_bram_5) and (not k12_needs_bram_5) and (not k23_needs_bram_5) and (not k22_needs_bram_5) and (not k21_needs_bram_5) and (not k20_needs_bram_5)));
	bram_12_input_sel(2) <= not ((k0_needs_bram_6 or k1_needs_bram_6 or k2_needs_bram_6 or k3_needs_bram_6) or ((k8_needs_bram_6 or k9_needs_bram_6 or k10_needs_bram_6 or k11_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k5_needs_bram_6) and (not k4_needs_bram_6)) or ((k16_needs_bram_6 or k17_needs_bram_6 or k18_needs_bram_6 or k19_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k5_needs_bram_6) and (not k4_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6) and (not k13_needs_bram_6) and (not k12_needs_bram_6)) or ((k24_needs_bram_6 or k25_needs_bram_6 or k26_needs_bram_6 or k27_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k5_needs_bram_6) and (not k4_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6) and (not k13_needs_bram_6) and (not k12_needs_bram_6) and (not k23_needs_bram_6) and (not k22_needs_bram_6) and (not k21_needs_bram_6) and (not k20_needs_bram_6)));
	bram_14_input_sel(2) <= not ((k0_needs_bram_7 or k1_needs_bram_7 or k2_needs_bram_7 or k3_needs_bram_7) or ((k8_needs_bram_7 or k9_needs_bram_7 or k10_needs_bram_7 or k11_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k5_needs_bram_7) and (not k4_needs_bram_7)) or ((k16_needs_bram_7 or k17_needs_bram_7 or k18_needs_bram_7 or k19_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k5_needs_bram_7) and (not k4_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7) and (not k13_needs_bram_7) and (not k12_needs_bram_7)) or ((k24_needs_bram_7 or k25_needs_bram_7 or k26_needs_bram_7 or k27_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k5_needs_bram_7) and (not k4_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7) and (not k13_needs_bram_7) and (not k12_needs_bram_7) and (not k23_needs_bram_7) and (not k22_needs_bram_7) and (not k21_needs_bram_7) and (not k20_needs_bram_7)));
	bram_16_input_sel(2) <= not ((k0_needs_bram_8 or k1_needs_bram_8 or k2_needs_bram_8 or k3_needs_bram_8) or ((k8_needs_bram_8 or k9_needs_bram_8 or k10_needs_bram_8 or k11_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k5_needs_bram_8) and (not k4_needs_bram_8)) or ((k16_needs_bram_8 or k17_needs_bram_8 or k18_needs_bram_8 or k19_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k5_needs_bram_8) and (not k4_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8) and (not k13_needs_bram_8) and (not k12_needs_bram_8)) or ((k24_needs_bram_8 or k25_needs_bram_8 or k26_needs_bram_8 or k27_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k5_needs_bram_8) and (not k4_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8) and (not k13_needs_bram_8) and (not k12_needs_bram_8) and (not k23_needs_bram_8) and (not k22_needs_bram_8) and (not k21_needs_bram_8) and (not k20_needs_bram_8)));
	bram_18_input_sel(2) <= not ((k0_needs_bram_9 or k1_needs_bram_9 or k2_needs_bram_9 or k3_needs_bram_9) or ((k8_needs_bram_9 or k9_needs_bram_9 or k10_needs_bram_9 or k11_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k5_needs_bram_9) and (not k4_needs_bram_9)) or ((k16_needs_bram_9 or k17_needs_bram_9 or k18_needs_bram_9 or k19_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k5_needs_bram_9) and (not k4_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9) and (not k13_needs_bram_9) and (not k12_needs_bram_9)) or ((k24_needs_bram_9 or k25_needs_bram_9 or k26_needs_bram_9 or k27_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k5_needs_bram_9) and (not k4_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9) and (not k13_needs_bram_9) and (not k12_needs_bram_9) and (not k23_needs_bram_9) and (not k22_needs_bram_9) and (not k21_needs_bram_9) and (not k20_needs_bram_9)));
	bram_20_input_sel(2) <= not ((k0_needs_bram_10 or k1_needs_bram_10 or k2_needs_bram_10 or k3_needs_bram_10) or ((k8_needs_bram_10 or k9_needs_bram_10 or k10_needs_bram_10 or k11_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k5_needs_bram_10) and (not k4_needs_bram_10)) or ((k16_needs_bram_10 or k17_needs_bram_10 or k18_needs_bram_10 or k19_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k5_needs_bram_10) and (not k4_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10) and (not k13_needs_bram_10) and (not k12_needs_bram_10)) or ((k24_needs_bram_10 or k25_needs_bram_10 or k26_needs_bram_10 or k27_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k5_needs_bram_10) and (not k4_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10) and (not k13_needs_bram_10) and (not k12_needs_bram_10) and (not k23_needs_bram_10) and (not k22_needs_bram_10) and (not k21_needs_bram_10) and (not k20_needs_bram_10)));
	bram_22_input_sel(2) <= not ((k0_needs_bram_11 or k1_needs_bram_11 or k2_needs_bram_11 or k3_needs_bram_11) or ((k8_needs_bram_11 or k9_needs_bram_11 or k10_needs_bram_11 or k11_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k5_needs_bram_11) and (not k4_needs_bram_11)) or ((k16_needs_bram_11 or k17_needs_bram_11 or k18_needs_bram_11 or k19_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k5_needs_bram_11) and (not k4_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11) and (not k13_needs_bram_11) and (not k12_needs_bram_11)) or ((k24_needs_bram_11 or k25_needs_bram_11 or k26_needs_bram_11 or k27_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k5_needs_bram_11) and (not k4_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11) and (not k13_needs_bram_11) and (not k12_needs_bram_11) and (not k23_needs_bram_11) and (not k22_needs_bram_11) and (not k21_needs_bram_11) and (not k20_needs_bram_11)));
	bram_24_input_sel(2) <= not ((k0_needs_bram_12 or k1_needs_bram_12 or k2_needs_bram_12 or k3_needs_bram_12) or ((k8_needs_bram_12 or k9_needs_bram_12 or k10_needs_bram_12 or k11_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k5_needs_bram_12) and (not k4_needs_bram_12)) or ((k16_needs_bram_12 or k17_needs_bram_12 or k18_needs_bram_12 or k19_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k5_needs_bram_12) and (not k4_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12) and (not k13_needs_bram_12) and (not k12_needs_bram_12)) or ((k24_needs_bram_12 or k25_needs_bram_12 or k26_needs_bram_12 or k27_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k5_needs_bram_12) and (not k4_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12) and (not k13_needs_bram_12) and (not k12_needs_bram_12) and (not k23_needs_bram_12) and (not k22_needs_bram_12) and (not k21_needs_bram_12) and (not k20_needs_bram_12)));
	bram_26_input_sel(2) <= not ((k0_needs_bram_13 or k1_needs_bram_13 or k2_needs_bram_13 or k3_needs_bram_13) or ((k8_needs_bram_13 or k9_needs_bram_13 or k10_needs_bram_13 or k11_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k5_needs_bram_13) and (not k4_needs_bram_13)) or ((k16_needs_bram_13 or k17_needs_bram_13 or k18_needs_bram_13 or k19_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k5_needs_bram_13) and (not k4_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13) and (not k13_needs_bram_13) and (not k12_needs_bram_13)) or ((k24_needs_bram_13 or k25_needs_bram_13 or k26_needs_bram_13 or k27_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k5_needs_bram_13) and (not k4_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13) and (not k13_needs_bram_13) and (not k12_needs_bram_13) and (not k23_needs_bram_13) and (not k22_needs_bram_13) and (not k21_needs_bram_13) and (not k20_needs_bram_13)));
	bram_28_input_sel(2) <= not ((k0_needs_bram_14 or k1_needs_bram_14 or k2_needs_bram_14 or k3_needs_bram_14) or ((k8_needs_bram_14 or k9_needs_bram_14 or k10_needs_bram_14 or k11_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k5_needs_bram_14) and (not k4_needs_bram_14)) or ((k16_needs_bram_14 or k17_needs_bram_14 or k18_needs_bram_14 or k19_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k5_needs_bram_14) and (not k4_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14) and (not k13_needs_bram_14) and (not k12_needs_bram_14)) or ((k24_needs_bram_14 or k25_needs_bram_14 or k26_needs_bram_14 or k27_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k5_needs_bram_14) and (not k4_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14) and (not k13_needs_bram_14) and (not k12_needs_bram_14) and (not k23_needs_bram_14) and (not k22_needs_bram_14) and (not k21_needs_bram_14) and (not k20_needs_bram_14)));
	bram_30_input_sel(2) <= not ((k0_needs_bram_15 or k1_needs_bram_15 or k2_needs_bram_15 or k3_needs_bram_15) or ((k8_needs_bram_15 or k9_needs_bram_15 or k10_needs_bram_15 or k11_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k5_needs_bram_15) and (not k4_needs_bram_15)) or ((k16_needs_bram_15 or k17_needs_bram_15 or k18_needs_bram_15 or k19_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k5_needs_bram_15) and (not k4_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15) and (not k13_needs_bram_15) and (not k12_needs_bram_15)) or ((k24_needs_bram_15 or k25_needs_bram_15 or k26_needs_bram_15 or k27_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k5_needs_bram_15) and (not k4_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15) and (not k13_needs_bram_15) and (not k12_needs_bram_15) and (not k23_needs_bram_15) and (not k22_needs_bram_15) and (not k21_needs_bram_15) and (not k20_needs_bram_15)));

	bram_0_input_sel(1) <= not ((k0_needs_bram_0 or k1_needs_bram_0) or ((k4_needs_bram_0 or k5_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0)) or ((k8_needs_bram_0 or k9_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0)) or ((k12_needs_bram_0 or k13_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k11_needs_bram_0) and (not k10_needs_bram_0)) or ((k16_needs_bram_0 or k17_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k11_needs_bram_0) and (not k10_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0)) or ((k20_needs_bram_0 or k21_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k11_needs_bram_0) and (not k10_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0) and (not k19_needs_bram_0) and (not k18_needs_bram_0)) or ((k24_needs_bram_0 or k25_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k11_needs_bram_0) and (not k10_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0) and (not k19_needs_bram_0) and (not k18_needs_bram_0) and (not k23_needs_bram_0) and (not k22_needs_bram_0)) or ((k28_needs_bram_0 or k29_needs_bram_0) and (not k3_needs_bram_0) and (not k2_needs_bram_0) and (not k7_needs_bram_0) and (not k6_needs_bram_0) and (not k11_needs_bram_0) and (not k10_needs_bram_0) and (not k15_needs_bram_0) and (not k14_needs_bram_0) and (not k19_needs_bram_0) and (not k18_needs_bram_0) and (not k23_needs_bram_0) and (not k22_needs_bram_0) and (not k27_needs_bram_0) and (not k26_needs_bram_0)));
	bram_2_input_sel(1) <= not ((k0_needs_bram_1 or k1_needs_bram_1) or ((k4_needs_bram_1 or k5_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1)) or ((k8_needs_bram_1 or k9_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1)) or ((k12_needs_bram_1 or k13_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k11_needs_bram_1) and (not k10_needs_bram_1)) or ((k16_needs_bram_1 or k17_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k11_needs_bram_1) and (not k10_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1)) or ((k20_needs_bram_1 or k21_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k11_needs_bram_1) and (not k10_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1) and (not k19_needs_bram_1) and (not k18_needs_bram_1)) or ((k24_needs_bram_1 or k25_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k11_needs_bram_1) and (not k10_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1) and (not k19_needs_bram_1) and (not k18_needs_bram_1) and (not k23_needs_bram_1) and (not k22_needs_bram_1)) or ((k28_needs_bram_1 or k29_needs_bram_1) and (not k3_needs_bram_1) and (not k2_needs_bram_1) and (not k7_needs_bram_1) and (not k6_needs_bram_1) and (not k11_needs_bram_1) and (not k10_needs_bram_1) and (not k15_needs_bram_1) and (not k14_needs_bram_1) and (not k19_needs_bram_1) and (not k18_needs_bram_1) and (not k23_needs_bram_1) and (not k22_needs_bram_1) and (not k27_needs_bram_1) and (not k26_needs_bram_1)));
	bram_4_input_sel(1) <= not ((k0_needs_bram_2 or k1_needs_bram_2) or ((k4_needs_bram_2 or k5_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2)) or ((k8_needs_bram_2 or k9_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2)) or ((k12_needs_bram_2 or k13_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k11_needs_bram_2) and (not k10_needs_bram_2)) or ((k16_needs_bram_2 or k17_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k11_needs_bram_2) and (not k10_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2)) or ((k20_needs_bram_2 or k21_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k11_needs_bram_2) and (not k10_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2) and (not k19_needs_bram_2) and (not k18_needs_bram_2)) or ((k24_needs_bram_2 or k25_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k11_needs_bram_2) and (not k10_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2) and (not k19_needs_bram_2) and (not k18_needs_bram_2) and (not k23_needs_bram_2) and (not k22_needs_bram_2)) or ((k28_needs_bram_2 or k29_needs_bram_2) and (not k3_needs_bram_2) and (not k2_needs_bram_2) and (not k7_needs_bram_2) and (not k6_needs_bram_2) and (not k11_needs_bram_2) and (not k10_needs_bram_2) and (not k15_needs_bram_2) and (not k14_needs_bram_2) and (not k19_needs_bram_2) and (not k18_needs_bram_2) and (not k23_needs_bram_2) and (not k22_needs_bram_2) and (not k27_needs_bram_2) and (not k26_needs_bram_2)));
	bram_6_input_sel(1) <= not ((k0_needs_bram_3 or k1_needs_bram_3) or ((k4_needs_bram_3 or k5_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3)) or ((k8_needs_bram_3 or k9_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3)) or ((k12_needs_bram_3 or k13_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k11_needs_bram_3) and (not k10_needs_bram_3)) or ((k16_needs_bram_3 or k17_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k11_needs_bram_3) and (not k10_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3)) or ((k20_needs_bram_3 or k21_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k11_needs_bram_3) and (not k10_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3) and (not k19_needs_bram_3) and (not k18_needs_bram_3)) or ((k24_needs_bram_3 or k25_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k11_needs_bram_3) and (not k10_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3) and (not k19_needs_bram_3) and (not k18_needs_bram_3) and (not k23_needs_bram_3) and (not k22_needs_bram_3)) or ((k28_needs_bram_3 or k29_needs_bram_3) and (not k3_needs_bram_3) and (not k2_needs_bram_3) and (not k7_needs_bram_3) and (not k6_needs_bram_3) and (not k11_needs_bram_3) and (not k10_needs_bram_3) and (not k15_needs_bram_3) and (not k14_needs_bram_3) and (not k19_needs_bram_3) and (not k18_needs_bram_3) and (not k23_needs_bram_3) and (not k22_needs_bram_3) and (not k27_needs_bram_3) and (not k26_needs_bram_3)));
	bram_8_input_sel(1) <= not ((k0_needs_bram_4 or k1_needs_bram_4) or ((k4_needs_bram_4 or k5_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4)) or ((k8_needs_bram_4 or k9_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4)) or ((k12_needs_bram_4 or k13_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k11_needs_bram_4) and (not k10_needs_bram_4)) or ((k16_needs_bram_4 or k17_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k11_needs_bram_4) and (not k10_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4)) or ((k20_needs_bram_4 or k21_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k11_needs_bram_4) and (not k10_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4) and (not k19_needs_bram_4) and (not k18_needs_bram_4)) or ((k24_needs_bram_4 or k25_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k11_needs_bram_4) and (not k10_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4) and (not k19_needs_bram_4) and (not k18_needs_bram_4) and (not k23_needs_bram_4) and (not k22_needs_bram_4)) or ((k28_needs_bram_4 or k29_needs_bram_4) and (not k3_needs_bram_4) and (not k2_needs_bram_4) and (not k7_needs_bram_4) and (not k6_needs_bram_4) and (not k11_needs_bram_4) and (not k10_needs_bram_4) and (not k15_needs_bram_4) and (not k14_needs_bram_4) and (not k19_needs_bram_4) and (not k18_needs_bram_4) and (not k23_needs_bram_4) and (not k22_needs_bram_4) and (not k27_needs_bram_4) and (not k26_needs_bram_4)));
	bram_10_input_sel(1) <= not ((k0_needs_bram_5 or k1_needs_bram_5) or ((k4_needs_bram_5 or k5_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5)) or ((k8_needs_bram_5 or k9_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5)) or ((k12_needs_bram_5 or k13_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k11_needs_bram_5) and (not k10_needs_bram_5)) or ((k16_needs_bram_5 or k17_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k11_needs_bram_5) and (not k10_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5)) or ((k20_needs_bram_5 or k21_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k11_needs_bram_5) and (not k10_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5) and (not k19_needs_bram_5) and (not k18_needs_bram_5)) or ((k24_needs_bram_5 or k25_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k11_needs_bram_5) and (not k10_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5) and (not k19_needs_bram_5) and (not k18_needs_bram_5) and (not k23_needs_bram_5) and (not k22_needs_bram_5)) or ((k28_needs_bram_5 or k29_needs_bram_5) and (not k3_needs_bram_5) and (not k2_needs_bram_5) and (not k7_needs_bram_5) and (not k6_needs_bram_5) and (not k11_needs_bram_5) and (not k10_needs_bram_5) and (not k15_needs_bram_5) and (not k14_needs_bram_5) and (not k19_needs_bram_5) and (not k18_needs_bram_5) and (not k23_needs_bram_5) and (not k22_needs_bram_5) and (not k27_needs_bram_5) and (not k26_needs_bram_5)));
	bram_12_input_sel(1) <= not ((k0_needs_bram_6 or k1_needs_bram_6) or ((k4_needs_bram_6 or k5_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6)) or ((k8_needs_bram_6 or k9_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6)) or ((k12_needs_bram_6 or k13_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k11_needs_bram_6) and (not k10_needs_bram_6)) or ((k16_needs_bram_6 or k17_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k11_needs_bram_6) and (not k10_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6)) or ((k20_needs_bram_6 or k21_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k11_needs_bram_6) and (not k10_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6) and (not k19_needs_bram_6) and (not k18_needs_bram_6)) or ((k24_needs_bram_6 or k25_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k11_needs_bram_6) and (not k10_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6) and (not k19_needs_bram_6) and (not k18_needs_bram_6) and (not k23_needs_bram_6) and (not k22_needs_bram_6)) or ((k28_needs_bram_6 or k29_needs_bram_6) and (not k3_needs_bram_6) and (not k2_needs_bram_6) and (not k7_needs_bram_6) and (not k6_needs_bram_6) and (not k11_needs_bram_6) and (not k10_needs_bram_6) and (not k15_needs_bram_6) and (not k14_needs_bram_6) and (not k19_needs_bram_6) and (not k18_needs_bram_6) and (not k23_needs_bram_6) and (not k22_needs_bram_6) and (not k27_needs_bram_6) and (not k26_needs_bram_6)));
	bram_14_input_sel(1) <= not ((k0_needs_bram_7 or k1_needs_bram_7) or ((k4_needs_bram_7 or k5_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7)) or ((k8_needs_bram_7 or k9_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7)) or ((k12_needs_bram_7 or k13_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k11_needs_bram_7) and (not k10_needs_bram_7)) or ((k16_needs_bram_7 or k17_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k11_needs_bram_7) and (not k10_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7)) or ((k20_needs_bram_7 or k21_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k11_needs_bram_7) and (not k10_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7) and (not k19_needs_bram_7) and (not k18_needs_bram_7)) or ((k24_needs_bram_7 or k25_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k11_needs_bram_7) and (not k10_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7) and (not k19_needs_bram_7) and (not k18_needs_bram_7) and (not k23_needs_bram_7) and (not k22_needs_bram_7)) or ((k28_needs_bram_7 or k29_needs_bram_7) and (not k3_needs_bram_7) and (not k2_needs_bram_7) and (not k7_needs_bram_7) and (not k6_needs_bram_7) and (not k11_needs_bram_7) and (not k10_needs_bram_7) and (not k15_needs_bram_7) and (not k14_needs_bram_7) and (not k19_needs_bram_7) and (not k18_needs_bram_7) and (not k23_needs_bram_7) and (not k22_needs_bram_7) and (not k27_needs_bram_7) and (not k26_needs_bram_7)));
	bram_16_input_sel(1) <= not ((k0_needs_bram_8 or k1_needs_bram_8) or ((k4_needs_bram_8 or k5_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8)) or ((k8_needs_bram_8 or k9_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8)) or ((k12_needs_bram_8 or k13_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k11_needs_bram_8) and (not k10_needs_bram_8)) or ((k16_needs_bram_8 or k17_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k11_needs_bram_8) and (not k10_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8)) or ((k20_needs_bram_8 or k21_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k11_needs_bram_8) and (not k10_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8) and (not k19_needs_bram_8) and (not k18_needs_bram_8)) or ((k24_needs_bram_8 or k25_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k11_needs_bram_8) and (not k10_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8) and (not k19_needs_bram_8) and (not k18_needs_bram_8) and (not k23_needs_bram_8) and (not k22_needs_bram_8)) or ((k28_needs_bram_8 or k29_needs_bram_8) and (not k3_needs_bram_8) and (not k2_needs_bram_8) and (not k7_needs_bram_8) and (not k6_needs_bram_8) and (not k11_needs_bram_8) and (not k10_needs_bram_8) and (not k15_needs_bram_8) and (not k14_needs_bram_8) and (not k19_needs_bram_8) and (not k18_needs_bram_8) and (not k23_needs_bram_8) and (not k22_needs_bram_8) and (not k27_needs_bram_8) and (not k26_needs_bram_8)));
	bram_18_input_sel(1) <= not ((k0_needs_bram_9 or k1_needs_bram_9) or ((k4_needs_bram_9 or k5_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9)) or ((k8_needs_bram_9 or k9_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9)) or ((k12_needs_bram_9 or k13_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k11_needs_bram_9) and (not k10_needs_bram_9)) or ((k16_needs_bram_9 or k17_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k11_needs_bram_9) and (not k10_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9)) or ((k20_needs_bram_9 or k21_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k11_needs_bram_9) and (not k10_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9) and (not k19_needs_bram_9) and (not k18_needs_bram_9)) or ((k24_needs_bram_9 or k25_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k11_needs_bram_9) and (not k10_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9) and (not k19_needs_bram_9) and (not k18_needs_bram_9) and (not k23_needs_bram_9) and (not k22_needs_bram_9)) or ((k28_needs_bram_9 or k29_needs_bram_9) and (not k3_needs_bram_9) and (not k2_needs_bram_9) and (not k7_needs_bram_9) and (not k6_needs_bram_9) and (not k11_needs_bram_9) and (not k10_needs_bram_9) and (not k15_needs_bram_9) and (not k14_needs_bram_9) and (not k19_needs_bram_9) and (not k18_needs_bram_9) and (not k23_needs_bram_9) and (not k22_needs_bram_9) and (not k27_needs_bram_9) and (not k26_needs_bram_9)));
	bram_20_input_sel(1) <= not ((k0_needs_bram_10 or k1_needs_bram_10) or ((k4_needs_bram_10 or k5_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10)) or ((k8_needs_bram_10 or k9_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10)) or ((k12_needs_bram_10 or k13_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k11_needs_bram_10) and (not k10_needs_bram_10)) or ((k16_needs_bram_10 or k17_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k11_needs_bram_10) and (not k10_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10)) or ((k20_needs_bram_10 or k21_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k11_needs_bram_10) and (not k10_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10) and (not k19_needs_bram_10) and (not k18_needs_bram_10)) or ((k24_needs_bram_10 or k25_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k11_needs_bram_10) and (not k10_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10) and (not k19_needs_bram_10) and (not k18_needs_bram_10) and (not k23_needs_bram_10) and (not k22_needs_bram_10)) or ((k28_needs_bram_10 or k29_needs_bram_10) and (not k3_needs_bram_10) and (not k2_needs_bram_10) and (not k7_needs_bram_10) and (not k6_needs_bram_10) and (not k11_needs_bram_10) and (not k10_needs_bram_10) and (not k15_needs_bram_10) and (not k14_needs_bram_10) and (not k19_needs_bram_10) and (not k18_needs_bram_10) and (not k23_needs_bram_10) and (not k22_needs_bram_10) and (not k27_needs_bram_10) and (not k26_needs_bram_10)));
	bram_22_input_sel(1) <= not ((k0_needs_bram_11 or k1_needs_bram_11) or ((k4_needs_bram_11 or k5_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11)) or ((k8_needs_bram_11 or k9_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11)) or ((k12_needs_bram_11 or k13_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k11_needs_bram_11) and (not k10_needs_bram_11)) or ((k16_needs_bram_11 or k17_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k11_needs_bram_11) and (not k10_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11)) or ((k20_needs_bram_11 or k21_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k11_needs_bram_11) and (not k10_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11) and (not k19_needs_bram_11) and (not k18_needs_bram_11)) or ((k24_needs_bram_11 or k25_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k11_needs_bram_11) and (not k10_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11) and (not k19_needs_bram_11) and (not k18_needs_bram_11) and (not k23_needs_bram_11) and (not k22_needs_bram_11)) or ((k28_needs_bram_11 or k29_needs_bram_11) and (not k3_needs_bram_11) and (not k2_needs_bram_11) and (not k7_needs_bram_11) and (not k6_needs_bram_11) and (not k11_needs_bram_11) and (not k10_needs_bram_11) and (not k15_needs_bram_11) and (not k14_needs_bram_11) and (not k19_needs_bram_11) and (not k18_needs_bram_11) and (not k23_needs_bram_11) and (not k22_needs_bram_11) and (not k27_needs_bram_11) and (not k26_needs_bram_11)));
	bram_24_input_sel(1) <= not ((k0_needs_bram_12 or k1_needs_bram_12) or ((k4_needs_bram_12 or k5_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12)) or ((k8_needs_bram_12 or k9_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12)) or ((k12_needs_bram_12 or k13_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k11_needs_bram_12) and (not k10_needs_bram_12)) or ((k16_needs_bram_12 or k17_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k11_needs_bram_12) and (not k10_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12)) or ((k20_needs_bram_12 or k21_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k11_needs_bram_12) and (not k10_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12) and (not k19_needs_bram_12) and (not k18_needs_bram_12)) or ((k24_needs_bram_12 or k25_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k11_needs_bram_12) and (not k10_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12) and (not k19_needs_bram_12) and (not k18_needs_bram_12) and (not k23_needs_bram_12) and (not k22_needs_bram_12)) or ((k28_needs_bram_12 or k29_needs_bram_12) and (not k3_needs_bram_12) and (not k2_needs_bram_12) and (not k7_needs_bram_12) and (not k6_needs_bram_12) and (not k11_needs_bram_12) and (not k10_needs_bram_12) and (not k15_needs_bram_12) and (not k14_needs_bram_12) and (not k19_needs_bram_12) and (not k18_needs_bram_12) and (not k23_needs_bram_12) and (not k22_needs_bram_12) and (not k27_needs_bram_12) and (not k26_needs_bram_12)));
	bram_26_input_sel(1) <= not ((k0_needs_bram_13 or k1_needs_bram_13) or ((k4_needs_bram_13 or k5_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13)) or ((k8_needs_bram_13 or k9_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13)) or ((k12_needs_bram_13 or k13_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k11_needs_bram_13) and (not k10_needs_bram_13)) or ((k16_needs_bram_13 or k17_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k11_needs_bram_13) and (not k10_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13)) or ((k20_needs_bram_13 or k21_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k11_needs_bram_13) and (not k10_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13) and (not k19_needs_bram_13) and (not k18_needs_bram_13)) or ((k24_needs_bram_13 or k25_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k11_needs_bram_13) and (not k10_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13) and (not k19_needs_bram_13) and (not k18_needs_bram_13) and (not k23_needs_bram_13) and (not k22_needs_bram_13)) or ((k28_needs_bram_13 or k29_needs_bram_13) and (not k3_needs_bram_13) and (not k2_needs_bram_13) and (not k7_needs_bram_13) and (not k6_needs_bram_13) and (not k11_needs_bram_13) and (not k10_needs_bram_13) and (not k15_needs_bram_13) and (not k14_needs_bram_13) and (not k19_needs_bram_13) and (not k18_needs_bram_13) and (not k23_needs_bram_13) and (not k22_needs_bram_13) and (not k27_needs_bram_13) and (not k26_needs_bram_13)));
	bram_28_input_sel(1) <= not ((k0_needs_bram_14 or k1_needs_bram_14) or ((k4_needs_bram_14 or k5_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14)) or ((k8_needs_bram_14 or k9_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14)) or ((k12_needs_bram_14 or k13_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k11_needs_bram_14) and (not k10_needs_bram_14)) or ((k16_needs_bram_14 or k17_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k11_needs_bram_14) and (not k10_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14)) or ((k20_needs_bram_14 or k21_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k11_needs_bram_14) and (not k10_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14) and (not k19_needs_bram_14) and (not k18_needs_bram_14)) or ((k24_needs_bram_14 or k25_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k11_needs_bram_14) and (not k10_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14) and (not k19_needs_bram_14) and (not k18_needs_bram_14) and (not k23_needs_bram_14) and (not k22_needs_bram_14)) or ((k28_needs_bram_14 or k29_needs_bram_14) and (not k3_needs_bram_14) and (not k2_needs_bram_14) and (not k7_needs_bram_14) and (not k6_needs_bram_14) and (not k11_needs_bram_14) and (not k10_needs_bram_14) and (not k15_needs_bram_14) and (not k14_needs_bram_14) and (not k19_needs_bram_14) and (not k18_needs_bram_14) and (not k23_needs_bram_14) and (not k22_needs_bram_14) and (not k27_needs_bram_14) and (not k26_needs_bram_14)));
	bram_30_input_sel(1) <= not ((k0_needs_bram_15 or k1_needs_bram_15) or ((k4_needs_bram_15 or k5_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15)) or ((k8_needs_bram_15 or k9_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15)) or ((k12_needs_bram_15 or k13_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k11_needs_bram_15) and (not k10_needs_bram_15)) or ((k16_needs_bram_15 or k17_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k11_needs_bram_15) and (not k10_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15)) or ((k20_needs_bram_15 or k21_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k11_needs_bram_15) and (not k10_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15) and (not k19_needs_bram_15) and (not k18_needs_bram_15)) or ((k24_needs_bram_15 or k25_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k11_needs_bram_15) and (not k10_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15) and (not k19_needs_bram_15) and (not k18_needs_bram_15) and (not k23_needs_bram_15) and (not k22_needs_bram_15)) or ((k28_needs_bram_15 or k29_needs_bram_15) and (not k3_needs_bram_15) and (not k2_needs_bram_15) and (not k7_needs_bram_15) and (not k6_needs_bram_15) and (not k11_needs_bram_15) and (not k10_needs_bram_15) and (not k15_needs_bram_15) and (not k14_needs_bram_15) and (not k19_needs_bram_15) and (not k18_needs_bram_15) and (not k23_needs_bram_15) and (not k22_needs_bram_15) and (not k27_needs_bram_15) and (not k26_needs_bram_15)));

	bram_0_input_sel(0) <= not ((k0_needs_bram_0) or ((k2_needs_bram_0) and (not k1_needs_bram_0)) or ((k4_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0)) or ((k6_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0)) or ((k8_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0)) or ((k10_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0)) or ((k12_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0)) or ((k14_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0)) or ((k16_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0)) or ((k18_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0)) or ((k20_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0) and (not k19_needs_bram_0)) or ((k22_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0) and (not k19_needs_bram_0) and (not k21_needs_bram_0)) or ((k24_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0) and (not k19_needs_bram_0) and (not k21_needs_bram_0) and (not k23_needs_bram_0)) or ((k26_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0) and (not k19_needs_bram_0) and (not k21_needs_bram_0) and (not k23_needs_bram_0) and (not k25_needs_bram_0)) or ((k28_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0) and (not k19_needs_bram_0) and (not k21_needs_bram_0) and (not k23_needs_bram_0) and (not k25_needs_bram_0) and (not k27_needs_bram_0)) or ((k30_needs_bram_0) and (not k1_needs_bram_0) and (not k3_needs_bram_0) and (not k5_needs_bram_0) and (not k7_needs_bram_0) and (not k9_needs_bram_0) and (not k11_needs_bram_0) and (not k13_needs_bram_0) and (not k15_needs_bram_0) and (not k17_needs_bram_0) and (not k19_needs_bram_0) and (not k21_needs_bram_0) and (not k23_needs_bram_0) and (not k25_needs_bram_0) and (not k27_needs_bram_0) and (not k29_needs_bram_0)));
	bram_2_input_sel(0) <= not ((k0_needs_bram_1) or ((k2_needs_bram_1) and (not k1_needs_bram_1)) or ((k4_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1)) or ((k6_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1)) or ((k8_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1)) or ((k10_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1)) or ((k12_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1)) or ((k14_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1)) or ((k16_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1)) or ((k18_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1)) or ((k20_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1) and (not k19_needs_bram_1)) or ((k22_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1) and (not k19_needs_bram_1) and (not k21_needs_bram_1)) or ((k24_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1) and (not k19_needs_bram_1) and (not k21_needs_bram_1) and (not k23_needs_bram_1)) or ((k26_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1) and (not k19_needs_bram_1) and (not k21_needs_bram_1) and (not k23_needs_bram_1) and (not k25_needs_bram_1)) or ((k28_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1) and (not k19_needs_bram_1) and (not k21_needs_bram_1) and (not k23_needs_bram_1) and (not k25_needs_bram_1) and (not k27_needs_bram_1)) or ((k30_needs_bram_1) and (not k1_needs_bram_1) and (not k3_needs_bram_1) and (not k5_needs_bram_1) and (not k7_needs_bram_1) and (not k9_needs_bram_1) and (not k11_needs_bram_1) and (not k13_needs_bram_1) and (not k15_needs_bram_1) and (not k17_needs_bram_1) and (not k19_needs_bram_1) and (not k21_needs_bram_1) and (not k23_needs_bram_1) and (not k25_needs_bram_1) and (not k27_needs_bram_1) and (not k29_needs_bram_1)));
	bram_4_input_sel(0) <= not ((k0_needs_bram_2) or ((k2_needs_bram_2) and (not k1_needs_bram_2)) or ((k4_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2)) or ((k6_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2)) or ((k8_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2)) or ((k10_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2)) or ((k12_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2)) or ((k14_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2)) or ((k16_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2)) or ((k18_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2)) or ((k20_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2) and (not k19_needs_bram_2)) or ((k22_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2) and (not k19_needs_bram_2) and (not k21_needs_bram_2)) or ((k24_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2) and (not k19_needs_bram_2) and (not k21_needs_bram_2) and (not k23_needs_bram_2)) or ((k26_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2) and (not k19_needs_bram_2) and (not k21_needs_bram_2) and (not k23_needs_bram_2) and (not k25_needs_bram_2)) or ((k28_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2) and (not k19_needs_bram_2) and (not k21_needs_bram_2) and (not k23_needs_bram_2) and (not k25_needs_bram_2) and (not k27_needs_bram_2)) or ((k30_needs_bram_2) and (not k1_needs_bram_2) and (not k3_needs_bram_2) and (not k5_needs_bram_2) and (not k7_needs_bram_2) and (not k9_needs_bram_2) and (not k11_needs_bram_2) and (not k13_needs_bram_2) and (not k15_needs_bram_2) and (not k17_needs_bram_2) and (not k19_needs_bram_2) and (not k21_needs_bram_2) and (not k23_needs_bram_2) and (not k25_needs_bram_2) and (not k27_needs_bram_2) and (not k29_needs_bram_2)));
	bram_6_input_sel(0) <= not ((k0_needs_bram_3) or ((k2_needs_bram_3) and (not k1_needs_bram_3)) or ((k4_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3)) or ((k6_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3)) or ((k8_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3)) or ((k10_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3)) or ((k12_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3)) or ((k14_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3)) or ((k16_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3)) or ((k18_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3)) or ((k20_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3) and (not k19_needs_bram_3)) or ((k22_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3) and (not k19_needs_bram_3) and (not k21_needs_bram_3)) or ((k24_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3) and (not k19_needs_bram_3) and (not k21_needs_bram_3) and (not k23_needs_bram_3)) or ((k26_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3) and (not k19_needs_bram_3) and (not k21_needs_bram_3) and (not k23_needs_bram_3) and (not k25_needs_bram_3)) or ((k28_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3) and (not k19_needs_bram_3) and (not k21_needs_bram_3) and (not k23_needs_bram_3) and (not k25_needs_bram_3) and (not k27_needs_bram_3)) or ((k30_needs_bram_3) and (not k1_needs_bram_3) and (not k3_needs_bram_3) and (not k5_needs_bram_3) and (not k7_needs_bram_3) and (not k9_needs_bram_3) and (not k11_needs_bram_3) and (not k13_needs_bram_3) and (not k15_needs_bram_3) and (not k17_needs_bram_3) and (not k19_needs_bram_3) and (not k21_needs_bram_3) and (not k23_needs_bram_3) and (not k25_needs_bram_3) and (not k27_needs_bram_3) and (not k29_needs_bram_3)));
	bram_8_input_sel(0) <= not ((k0_needs_bram_4) or ((k2_needs_bram_4) and (not k1_needs_bram_4)) or ((k4_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4)) or ((k6_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4)) or ((k8_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4)) or ((k10_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4)) or ((k12_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4)) or ((k14_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4)) or ((k16_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4)) or ((k18_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4)) or ((k20_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4) and (not k19_needs_bram_4)) or ((k22_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4) and (not k19_needs_bram_4) and (not k21_needs_bram_4)) or ((k24_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4) and (not k19_needs_bram_4) and (not k21_needs_bram_4) and (not k23_needs_bram_4)) or ((k26_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4) and (not k19_needs_bram_4) and (not k21_needs_bram_4) and (not k23_needs_bram_4) and (not k25_needs_bram_4)) or ((k28_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4) and (not k19_needs_bram_4) and (not k21_needs_bram_4) and (not k23_needs_bram_4) and (not k25_needs_bram_4) and (not k27_needs_bram_4)) or ((k30_needs_bram_4) and (not k1_needs_bram_4) and (not k3_needs_bram_4) and (not k5_needs_bram_4) and (not k7_needs_bram_4) and (not k9_needs_bram_4) and (not k11_needs_bram_4) and (not k13_needs_bram_4) and (not k15_needs_bram_4) and (not k17_needs_bram_4) and (not k19_needs_bram_4) and (not k21_needs_bram_4) and (not k23_needs_bram_4) and (not k25_needs_bram_4) and (not k27_needs_bram_4) and (not k29_needs_bram_4)));
	bram_10_input_sel(0) <= not ((k0_needs_bram_5) or ((k2_needs_bram_5) and (not k1_needs_bram_5)) or ((k4_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5)) or ((k6_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5)) or ((k8_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5)) or ((k10_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5)) or ((k12_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5)) or ((k14_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5)) or ((k16_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5)) or ((k18_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5)) or ((k20_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5) and (not k19_needs_bram_5)) or ((k22_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5) and (not k19_needs_bram_5) and (not k21_needs_bram_5)) or ((k24_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5) and (not k19_needs_bram_5) and (not k21_needs_bram_5) and (not k23_needs_bram_5)) or ((k26_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5) and (not k19_needs_bram_5) and (not k21_needs_bram_5) and (not k23_needs_bram_5) and (not k25_needs_bram_5)) or ((k28_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5) and (not k19_needs_bram_5) and (not k21_needs_bram_5) and (not k23_needs_bram_5) and (not k25_needs_bram_5) and (not k27_needs_bram_5)) or ((k30_needs_bram_5) and (not k1_needs_bram_5) and (not k3_needs_bram_5) and (not k5_needs_bram_5) and (not k7_needs_bram_5) and (not k9_needs_bram_5) and (not k11_needs_bram_5) and (not k13_needs_bram_5) and (not k15_needs_bram_5) and (not k17_needs_bram_5) and (not k19_needs_bram_5) and (not k21_needs_bram_5) and (not k23_needs_bram_5) and (not k25_needs_bram_5) and (not k27_needs_bram_5) and (not k29_needs_bram_5)));
	bram_12_input_sel(0) <= not ((k0_needs_bram_6) or ((k2_needs_bram_6) and (not k1_needs_bram_6)) or ((k4_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6)) or ((k6_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6)) or ((k8_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6)) or ((k10_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6)) or ((k12_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6)) or ((k14_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6)) or ((k16_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6)) or ((k18_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6)) or ((k20_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6) and (not k19_needs_bram_6)) or ((k22_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6) and (not k19_needs_bram_6) and (not k21_needs_bram_6)) or ((k24_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6) and (not k19_needs_bram_6) and (not k21_needs_bram_6) and (not k23_needs_bram_6)) or ((k26_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6) and (not k19_needs_bram_6) and (not k21_needs_bram_6) and (not k23_needs_bram_6) and (not k25_needs_bram_6)) or ((k28_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6) and (not k19_needs_bram_6) and (not k21_needs_bram_6) and (not k23_needs_bram_6) and (not k25_needs_bram_6) and (not k27_needs_bram_6)) or ((k30_needs_bram_6) and (not k1_needs_bram_6) and (not k3_needs_bram_6) and (not k5_needs_bram_6) and (not k7_needs_bram_6) and (not k9_needs_bram_6) and (not k11_needs_bram_6) and (not k13_needs_bram_6) and (not k15_needs_bram_6) and (not k17_needs_bram_6) and (not k19_needs_bram_6) and (not k21_needs_bram_6) and (not k23_needs_bram_6) and (not k25_needs_bram_6) and (not k27_needs_bram_6) and (not k29_needs_bram_6)));
	bram_14_input_sel(0) <= not ((k0_needs_bram_7) or ((k2_needs_bram_7) and (not k1_needs_bram_7)) or ((k4_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7)) or ((k6_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7)) or ((k8_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7)) or ((k10_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7)) or ((k12_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7)) or ((k14_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7)) or ((k16_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7)) or ((k18_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7)) or ((k20_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7) and (not k19_needs_bram_7)) or ((k22_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7) and (not k19_needs_bram_7) and (not k21_needs_bram_7)) or ((k24_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7) and (not k19_needs_bram_7) and (not k21_needs_bram_7) and (not k23_needs_bram_7)) or ((k26_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7) and (not k19_needs_bram_7) and (not k21_needs_bram_7) and (not k23_needs_bram_7) and (not k25_needs_bram_7)) or ((k28_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7) and (not k19_needs_bram_7) and (not k21_needs_bram_7) and (not k23_needs_bram_7) and (not k25_needs_bram_7) and (not k27_needs_bram_7)) or ((k30_needs_bram_7) and (not k1_needs_bram_7) and (not k3_needs_bram_7) and (not k5_needs_bram_7) and (not k7_needs_bram_7) and (not k9_needs_bram_7) and (not k11_needs_bram_7) and (not k13_needs_bram_7) and (not k15_needs_bram_7) and (not k17_needs_bram_7) and (not k19_needs_bram_7) and (not k21_needs_bram_7) and (not k23_needs_bram_7) and (not k25_needs_bram_7) and (not k27_needs_bram_7) and (not k29_needs_bram_7)));
	bram_16_input_sel(0) <= not ((k0_needs_bram_8) or ((k2_needs_bram_8) and (not k1_needs_bram_8)) or ((k4_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8)) or ((k6_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8)) or ((k8_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8)) or ((k10_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8)) or ((k12_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8)) or ((k14_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8)) or ((k16_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8)) or ((k18_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8)) or ((k20_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8) and (not k19_needs_bram_8)) or ((k22_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8) and (not k19_needs_bram_8) and (not k21_needs_bram_8)) or ((k24_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8) and (not k19_needs_bram_8) and (not k21_needs_bram_8) and (not k23_needs_bram_8)) or ((k26_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8) and (not k19_needs_bram_8) and (not k21_needs_bram_8) and (not k23_needs_bram_8) and (not k25_needs_bram_8)) or ((k28_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8) and (not k19_needs_bram_8) and (not k21_needs_bram_8) and (not k23_needs_bram_8) and (not k25_needs_bram_8) and (not k27_needs_bram_8)) or ((k30_needs_bram_8) and (not k1_needs_bram_8) and (not k3_needs_bram_8) and (not k5_needs_bram_8) and (not k7_needs_bram_8) and (not k9_needs_bram_8) and (not k11_needs_bram_8) and (not k13_needs_bram_8) and (not k15_needs_bram_8) and (not k17_needs_bram_8) and (not k19_needs_bram_8) and (not k21_needs_bram_8) and (not k23_needs_bram_8) and (not k25_needs_bram_8) and (not k27_needs_bram_8) and (not k29_needs_bram_8)));
	bram_18_input_sel(0) <= not ((k0_needs_bram_9) or ((k2_needs_bram_9) and (not k1_needs_bram_9)) or ((k4_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9)) or ((k6_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9)) or ((k8_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9)) or ((k10_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9)) or ((k12_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9)) or ((k14_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9)) or ((k16_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9)) or ((k18_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9)) or ((k20_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9) and (not k19_needs_bram_9)) or ((k22_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9) and (not k19_needs_bram_9) and (not k21_needs_bram_9)) or ((k24_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9) and (not k19_needs_bram_9) and (not k21_needs_bram_9) and (not k23_needs_bram_9)) or ((k26_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9) and (not k19_needs_bram_9) and (not k21_needs_bram_9) and (not k23_needs_bram_9) and (not k25_needs_bram_9)) or ((k28_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9) and (not k19_needs_bram_9) and (not k21_needs_bram_9) and (not k23_needs_bram_9) and (not k25_needs_bram_9) and (not k27_needs_bram_9)) or ((k30_needs_bram_9) and (not k1_needs_bram_9) and (not k3_needs_bram_9) and (not k5_needs_bram_9) and (not k7_needs_bram_9) and (not k9_needs_bram_9) and (not k11_needs_bram_9) and (not k13_needs_bram_9) and (not k15_needs_bram_9) and (not k17_needs_bram_9) and (not k19_needs_bram_9) and (not k21_needs_bram_9) and (not k23_needs_bram_9) and (not k25_needs_bram_9) and (not k27_needs_bram_9) and (not k29_needs_bram_9)));
	bram_20_input_sel(0) <= not ((k0_needs_bram_10) or ((k2_needs_bram_10) and (not k1_needs_bram_10)) or ((k4_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10)) or ((k6_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10)) or ((k8_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10)) or ((k10_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10)) or ((k12_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10)) or ((k14_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10)) or ((k16_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10)) or ((k18_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10)) or ((k20_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10) and (not k19_needs_bram_10)) or ((k22_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10) and (not k19_needs_bram_10) and (not k21_needs_bram_10)) or ((k24_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10) and (not k19_needs_bram_10) and (not k21_needs_bram_10) and (not k23_needs_bram_10)) or ((k26_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10) and (not k19_needs_bram_10) and (not k21_needs_bram_10) and (not k23_needs_bram_10) and (not k25_needs_bram_10)) or ((k28_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10) and (not k19_needs_bram_10) and (not k21_needs_bram_10) and (not k23_needs_bram_10) and (not k25_needs_bram_10) and (not k27_needs_bram_10)) or ((k30_needs_bram_10) and (not k1_needs_bram_10) and (not k3_needs_bram_10) and (not k5_needs_bram_10) and (not k7_needs_bram_10) and (not k9_needs_bram_10) and (not k11_needs_bram_10) and (not k13_needs_bram_10) and (not k15_needs_bram_10) and (not k17_needs_bram_10) and (not k19_needs_bram_10) and (not k21_needs_bram_10) and (not k23_needs_bram_10) and (not k25_needs_bram_10) and (not k27_needs_bram_10) and (not k29_needs_bram_10)));
	bram_22_input_sel(0) <= not ((k0_needs_bram_11) or ((k2_needs_bram_11) and (not k1_needs_bram_11)) or ((k4_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11)) or ((k6_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11)) or ((k8_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11)) or ((k10_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11)) or ((k12_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11)) or ((k14_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11)) or ((k16_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11)) or ((k18_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11)) or ((k20_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11) and (not k19_needs_bram_11)) or ((k22_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11) and (not k19_needs_bram_11) and (not k21_needs_bram_11)) or ((k24_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11) and (not k19_needs_bram_11) and (not k21_needs_bram_11) and (not k23_needs_bram_11)) or ((k26_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11) and (not k19_needs_bram_11) and (not k21_needs_bram_11) and (not k23_needs_bram_11) and (not k25_needs_bram_11)) or ((k28_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11) and (not k19_needs_bram_11) and (not k21_needs_bram_11) and (not k23_needs_bram_11) and (not k25_needs_bram_11) and (not k27_needs_bram_11)) or ((k30_needs_bram_11) and (not k1_needs_bram_11) and (not k3_needs_bram_11) and (not k5_needs_bram_11) and (not k7_needs_bram_11) and (not k9_needs_bram_11) and (not k11_needs_bram_11) and (not k13_needs_bram_11) and (not k15_needs_bram_11) and (not k17_needs_bram_11) and (not k19_needs_bram_11) and (not k21_needs_bram_11) and (not k23_needs_bram_11) and (not k25_needs_bram_11) and (not k27_needs_bram_11) and (not k29_needs_bram_11)));
	bram_24_input_sel(0) <= not ((k0_needs_bram_12) or ((k2_needs_bram_12) and (not k1_needs_bram_12)) or ((k4_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12)) or ((k6_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12)) or ((k8_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12)) or ((k10_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12)) or ((k12_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12)) or ((k14_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12)) or ((k16_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12)) or ((k18_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12)) or ((k20_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12) and (not k19_needs_bram_12)) or ((k22_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12) and (not k19_needs_bram_12) and (not k21_needs_bram_12)) or ((k24_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12) and (not k19_needs_bram_12) and (not k21_needs_bram_12) and (not k23_needs_bram_12)) or ((k26_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12) and (not k19_needs_bram_12) and (not k21_needs_bram_12) and (not k23_needs_bram_12) and (not k25_needs_bram_12)) or ((k28_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12) and (not k19_needs_bram_12) and (not k21_needs_bram_12) and (not k23_needs_bram_12) and (not k25_needs_bram_12) and (not k27_needs_bram_12)) or ((k30_needs_bram_12) and (not k1_needs_bram_12) and (not k3_needs_bram_12) and (not k5_needs_bram_12) and (not k7_needs_bram_12) and (not k9_needs_bram_12) and (not k11_needs_bram_12) and (not k13_needs_bram_12) and (not k15_needs_bram_12) and (not k17_needs_bram_12) and (not k19_needs_bram_12) and (not k21_needs_bram_12) and (not k23_needs_bram_12) and (not k25_needs_bram_12) and (not k27_needs_bram_12) and (not k29_needs_bram_12)));
	bram_26_input_sel(0) <= not ((k0_needs_bram_13) or ((k2_needs_bram_13) and (not k1_needs_bram_13)) or ((k4_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13)) or ((k6_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13)) or ((k8_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13)) or ((k10_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13)) or ((k12_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13)) or ((k14_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13)) or ((k16_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13)) or ((k18_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13)) or ((k20_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13) and (not k19_needs_bram_13)) or ((k22_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13) and (not k19_needs_bram_13) and (not k21_needs_bram_13)) or ((k24_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13) and (not k19_needs_bram_13) and (not k21_needs_bram_13) and (not k23_needs_bram_13)) or ((k26_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13) and (not k19_needs_bram_13) and (not k21_needs_bram_13) and (not k23_needs_bram_13) and (not k25_needs_bram_13)) or ((k28_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13) and (not k19_needs_bram_13) and (not k21_needs_bram_13) and (not k23_needs_bram_13) and (not k25_needs_bram_13) and (not k27_needs_bram_13)) or ((k30_needs_bram_13) and (not k1_needs_bram_13) and (not k3_needs_bram_13) and (not k5_needs_bram_13) and (not k7_needs_bram_13) and (not k9_needs_bram_13) and (not k11_needs_bram_13) and (not k13_needs_bram_13) and (not k15_needs_bram_13) and (not k17_needs_bram_13) and (not k19_needs_bram_13) and (not k21_needs_bram_13) and (not k23_needs_bram_13) and (not k25_needs_bram_13) and (not k27_needs_bram_13) and (not k29_needs_bram_13)));
	bram_28_input_sel(0) <= not ((k0_needs_bram_14) or ((k2_needs_bram_14) and (not k1_needs_bram_14)) or ((k4_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14)) or ((k6_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14)) or ((k8_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14)) or ((k10_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14)) or ((k12_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14)) or ((k14_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14)) or ((k16_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14)) or ((k18_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14)) or ((k20_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14) and (not k19_needs_bram_14)) or ((k22_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14) and (not k19_needs_bram_14) and (not k21_needs_bram_14)) or ((k24_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14) and (not k19_needs_bram_14) and (not k21_needs_bram_14) and (not k23_needs_bram_14)) or ((k26_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14) and (not k19_needs_bram_14) and (not k21_needs_bram_14) and (not k23_needs_bram_14) and (not k25_needs_bram_14)) or ((k28_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14) and (not k19_needs_bram_14) and (not k21_needs_bram_14) and (not k23_needs_bram_14) and (not k25_needs_bram_14) and (not k27_needs_bram_14)) or ((k30_needs_bram_14) and (not k1_needs_bram_14) and (not k3_needs_bram_14) and (not k5_needs_bram_14) and (not k7_needs_bram_14) and (not k9_needs_bram_14) and (not k11_needs_bram_14) and (not k13_needs_bram_14) and (not k15_needs_bram_14) and (not k17_needs_bram_14) and (not k19_needs_bram_14) and (not k21_needs_bram_14) and (not k23_needs_bram_14) and (not k25_needs_bram_14) and (not k27_needs_bram_14) and (not k29_needs_bram_14)));
	bram_30_input_sel(0) <= not ((k0_needs_bram_15) or ((k2_needs_bram_15) and (not k1_needs_bram_15)) or ((k4_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15)) or ((k6_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15)) or ((k8_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15)) or ((k10_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15)) or ((k12_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15)) or ((k14_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15)) or ((k16_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15)) or ((k18_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15)) or ((k20_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15) and (not k19_needs_bram_15)) or ((k22_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15) and (not k19_needs_bram_15) and (not k21_needs_bram_15)) or ((k24_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15) and (not k19_needs_bram_15) and (not k21_needs_bram_15) and (not k23_needs_bram_15)) or ((k26_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15) and (not k19_needs_bram_15) and (not k21_needs_bram_15) and (not k23_needs_bram_15) and (not k25_needs_bram_15)) or ((k28_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15) and (not k19_needs_bram_15) and (not k21_needs_bram_15) and (not k23_needs_bram_15) and (not k25_needs_bram_15) and (not k27_needs_bram_15)) or ((k30_needs_bram_15) and (not k1_needs_bram_15) and (not k3_needs_bram_15) and (not k5_needs_bram_15) and (not k7_needs_bram_15) and (not k9_needs_bram_15) and (not k11_needs_bram_15) and (not k13_needs_bram_15) and (not k15_needs_bram_15) and (not k17_needs_bram_15) and (not k19_needs_bram_15) and (not k21_needs_bram_15) and (not k23_needs_bram_15) and (not k25_needs_bram_15) and (not k27_needs_bram_15) and (not k29_needs_bram_15)));


	bram_1_input_sel(4) <= (k31_needs_bram_0 or k30_needs_bram_0 or k29_needs_bram_0 or k28_needs_bram_0 or k27_needs_bram_0 or k26_needs_bram_0 or k25_needs_bram_0 or k24_needs_bram_0 or k23_needs_bram_0 or k22_needs_bram_0 or k21_needs_bram_0 or k20_needs_bram_0 or k19_needs_bram_0 or k18_needs_bram_0 or k17_needs_bram_0 or k16_needs_bram_0);
	bram_3_input_sel(4) <= (k31_needs_bram_1 or k30_needs_bram_1 or k29_needs_bram_1 or k28_needs_bram_1 or k27_needs_bram_1 or k26_needs_bram_1 or k25_needs_bram_1 or k24_needs_bram_1 or k23_needs_bram_1 or k22_needs_bram_1 or k21_needs_bram_1 or k20_needs_bram_1 or k19_needs_bram_1 or k18_needs_bram_1 or k17_needs_bram_1 or k16_needs_bram_1);
	bram_5_input_sel(4) <= (k31_needs_bram_2 or k30_needs_bram_2 or k29_needs_bram_2 or k28_needs_bram_2 or k27_needs_bram_2 or k26_needs_bram_2 or k25_needs_bram_2 or k24_needs_bram_2 or k23_needs_bram_2 or k22_needs_bram_2 or k21_needs_bram_2 or k20_needs_bram_2 or k19_needs_bram_2 or k18_needs_bram_2 or k17_needs_bram_2 or k16_needs_bram_2);
	bram_7_input_sel(4) <= (k31_needs_bram_3 or k30_needs_bram_3 or k29_needs_bram_3 or k28_needs_bram_3 or k27_needs_bram_3 or k26_needs_bram_3 or k25_needs_bram_3 or k24_needs_bram_3 or k23_needs_bram_3 or k22_needs_bram_3 or k21_needs_bram_3 or k20_needs_bram_3 or k19_needs_bram_3 or k18_needs_bram_3 or k17_needs_bram_3 or k16_needs_bram_3);
	bram_9_input_sel(4) <= (k31_needs_bram_4 or k30_needs_bram_4 or k29_needs_bram_4 or k28_needs_bram_4 or k27_needs_bram_4 or k26_needs_bram_4 or k25_needs_bram_4 or k24_needs_bram_4 or k23_needs_bram_4 or k22_needs_bram_4 or k21_needs_bram_4 or k20_needs_bram_4 or k19_needs_bram_4 or k18_needs_bram_4 or k17_needs_bram_4 or k16_needs_bram_4);
	bram_11_input_sel(4) <= (k31_needs_bram_5 or k30_needs_bram_5 or k29_needs_bram_5 or k28_needs_bram_5 or k27_needs_bram_5 or k26_needs_bram_5 or k25_needs_bram_5 or k24_needs_bram_5 or k23_needs_bram_5 or k22_needs_bram_5 or k21_needs_bram_5 or k20_needs_bram_5 or k19_needs_bram_5 or k18_needs_bram_5 or k17_needs_bram_5 or k16_needs_bram_5);
	bram_13_input_sel(4) <= (k31_needs_bram_6 or k30_needs_bram_6 or k29_needs_bram_6 or k28_needs_bram_6 or k27_needs_bram_6 or k26_needs_bram_6 or k25_needs_bram_6 or k24_needs_bram_6 or k23_needs_bram_6 or k22_needs_bram_6 or k21_needs_bram_6 or k20_needs_bram_6 or k19_needs_bram_6 or k18_needs_bram_6 or k17_needs_bram_6 or k16_needs_bram_6);
	bram_15_input_sel(4) <= (k31_needs_bram_7 or k30_needs_bram_7 or k29_needs_bram_7 or k28_needs_bram_7 or k27_needs_bram_7 or k26_needs_bram_7 or k25_needs_bram_7 or k24_needs_bram_7 or k23_needs_bram_7 or k22_needs_bram_7 or k21_needs_bram_7 or k20_needs_bram_7 or k19_needs_bram_7 or k18_needs_bram_7 or k17_needs_bram_7 or k16_needs_bram_7);
	bram_17_input_sel(4) <= (k31_needs_bram_8 or k30_needs_bram_8 or k29_needs_bram_8 or k28_needs_bram_8 or k27_needs_bram_8 or k26_needs_bram_8 or k25_needs_bram_8 or k24_needs_bram_8 or k23_needs_bram_8 or k22_needs_bram_8 or k21_needs_bram_8 or k20_needs_bram_8 or k19_needs_bram_8 or k18_needs_bram_8 or k17_needs_bram_8 or k16_needs_bram_8);
	bram_19_input_sel(4) <= (k31_needs_bram_9 or k30_needs_bram_9 or k29_needs_bram_9 or k28_needs_bram_9 or k27_needs_bram_9 or k26_needs_bram_9 or k25_needs_bram_9 or k24_needs_bram_9 or k23_needs_bram_9 or k22_needs_bram_9 or k21_needs_bram_9 or k20_needs_bram_9 or k19_needs_bram_9 or k18_needs_bram_9 or k17_needs_bram_9 or k16_needs_bram_9);
	bram_21_input_sel(4) <= (k31_needs_bram_10 or k30_needs_bram_10 or k29_needs_bram_10 or k28_needs_bram_10 or k27_needs_bram_10 or k26_needs_bram_10 or k25_needs_bram_10 or k24_needs_bram_10 or k23_needs_bram_10 or k22_needs_bram_10 or k21_needs_bram_10 or k20_needs_bram_10 or k19_needs_bram_10 or k18_needs_bram_10 or k17_needs_bram_10 or k16_needs_bram_10);
	bram_23_input_sel(4) <= (k31_needs_bram_11 or k30_needs_bram_11 or k29_needs_bram_11 or k28_needs_bram_11 or k27_needs_bram_11 or k26_needs_bram_11 or k25_needs_bram_11 or k24_needs_bram_11 or k23_needs_bram_11 or k22_needs_bram_11 or k21_needs_bram_11 or k20_needs_bram_11 or k19_needs_bram_11 or k18_needs_bram_11 or k17_needs_bram_11 or k16_needs_bram_11);
	bram_25_input_sel(4) <= (k31_needs_bram_12 or k30_needs_bram_12 or k29_needs_bram_12 or k28_needs_bram_12 or k27_needs_bram_12 or k26_needs_bram_12 or k25_needs_bram_12 or k24_needs_bram_12 or k23_needs_bram_12 or k22_needs_bram_12 or k21_needs_bram_12 or k20_needs_bram_12 or k19_needs_bram_12 or k18_needs_bram_12 or k17_needs_bram_12 or k16_needs_bram_12);
	bram_27_input_sel(4) <= (k31_needs_bram_13 or k30_needs_bram_13 or k29_needs_bram_13 or k28_needs_bram_13 or k27_needs_bram_13 or k26_needs_bram_13 or k25_needs_bram_13 or k24_needs_bram_13 or k23_needs_bram_13 or k22_needs_bram_13 or k21_needs_bram_13 or k20_needs_bram_13 or k19_needs_bram_13 or k18_needs_bram_13 or k17_needs_bram_13 or k16_needs_bram_13);
	bram_29_input_sel(4) <= (k31_needs_bram_14 or k30_needs_bram_14 or k29_needs_bram_14 or k28_needs_bram_14 or k27_needs_bram_14 or k26_needs_bram_14 or k25_needs_bram_14 or k24_needs_bram_14 or k23_needs_bram_14 or k22_needs_bram_14 or k21_needs_bram_14 or k20_needs_bram_14 or k19_needs_bram_14 or k18_needs_bram_14 or k17_needs_bram_14 or k16_needs_bram_14);
	bram_31_input_sel(4) <= (k31_needs_bram_15 or k30_needs_bram_15 or k29_needs_bram_15 or k28_needs_bram_15 or k27_needs_bram_15 or k26_needs_bram_15 or k25_needs_bram_15 or k24_needs_bram_15 or k23_needs_bram_15 or k22_needs_bram_15 or k21_needs_bram_15 or k20_needs_bram_15 or k19_needs_bram_15 or k18_needs_bram_15 or k17_needs_bram_15 or k16_needs_bram_15);

	bram_1_input_sel(3) <= (k31_needs_bram_0 or k30_needs_bram_0 or k29_needs_bram_0 or k28_needs_bram_0 or k27_needs_bram_0 or k26_needs_bram_0 or k25_needs_bram_0 or k24_needs_bram_0) or ((k15_needs_bram_0 or k14_needs_bram_0 or k13_needs_bram_0 or k12_needs_bram_0 or k11_needs_bram_0 or k10_needs_bram_0 or k9_needs_bram_0 or k8_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0) and (not k18_needs_bram_0) and (not k19_needs_bram_0) and (not k20_needs_bram_0) and (not k21_needs_bram_0) and (not k22_needs_bram_0) and (not k23_needs_bram_0));
	bram_3_input_sel(3) <= (k31_needs_bram_1 or k30_needs_bram_1 or k29_needs_bram_1 or k28_needs_bram_1 or k27_needs_bram_1 or k26_needs_bram_1 or k25_needs_bram_1 or k24_needs_bram_1) or ((k15_needs_bram_1 or k14_needs_bram_1 or k13_needs_bram_1 or k12_needs_bram_1 or k11_needs_bram_1 or k10_needs_bram_1 or k9_needs_bram_1 or k8_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1) and (not k18_needs_bram_1) and (not k19_needs_bram_1) and (not k20_needs_bram_1) and (not k21_needs_bram_1) and (not k22_needs_bram_1) and (not k23_needs_bram_1));
	bram_5_input_sel(3) <= (k31_needs_bram_2 or k30_needs_bram_2 or k29_needs_bram_2 or k28_needs_bram_2 or k27_needs_bram_2 or k26_needs_bram_2 or k25_needs_bram_2 or k24_needs_bram_2) or ((k15_needs_bram_2 or k14_needs_bram_2 or k13_needs_bram_2 or k12_needs_bram_2 or k11_needs_bram_2 or k10_needs_bram_2 or k9_needs_bram_2 or k8_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2) and (not k18_needs_bram_2) and (not k19_needs_bram_2) and (not k20_needs_bram_2) and (not k21_needs_bram_2) and (not k22_needs_bram_2) and (not k23_needs_bram_2));
	bram_7_input_sel(3) <= (k31_needs_bram_3 or k30_needs_bram_3 or k29_needs_bram_3 or k28_needs_bram_3 or k27_needs_bram_3 or k26_needs_bram_3 or k25_needs_bram_3 or k24_needs_bram_3) or ((k15_needs_bram_3 or k14_needs_bram_3 or k13_needs_bram_3 or k12_needs_bram_3 or k11_needs_bram_3 or k10_needs_bram_3 or k9_needs_bram_3 or k8_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3) and (not k18_needs_bram_3) and (not k19_needs_bram_3) and (not k20_needs_bram_3) and (not k21_needs_bram_3) and (not k22_needs_bram_3) and (not k23_needs_bram_3));
	bram_9_input_sel(3) <= (k31_needs_bram_4 or k30_needs_bram_4 or k29_needs_bram_4 or k28_needs_bram_4 or k27_needs_bram_4 or k26_needs_bram_4 or k25_needs_bram_4 or k24_needs_bram_4) or ((k15_needs_bram_4 or k14_needs_bram_4 or k13_needs_bram_4 or k12_needs_bram_4 or k11_needs_bram_4 or k10_needs_bram_4 or k9_needs_bram_4 or k8_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4) and (not k18_needs_bram_4) and (not k19_needs_bram_4) and (not k20_needs_bram_4) and (not k21_needs_bram_4) and (not k22_needs_bram_4) and (not k23_needs_bram_4));
	bram_11_input_sel(3) <= (k31_needs_bram_5 or k30_needs_bram_5 or k29_needs_bram_5 or k28_needs_bram_5 or k27_needs_bram_5 or k26_needs_bram_5 or k25_needs_bram_5 or k24_needs_bram_5) or ((k15_needs_bram_5 or k14_needs_bram_5 or k13_needs_bram_5 or k12_needs_bram_5 or k11_needs_bram_5 or k10_needs_bram_5 or k9_needs_bram_5 or k8_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5) and (not k18_needs_bram_5) and (not k19_needs_bram_5) and (not k20_needs_bram_5) and (not k21_needs_bram_5) and (not k22_needs_bram_5) and (not k23_needs_bram_5));
	bram_13_input_sel(3) <= (k31_needs_bram_6 or k30_needs_bram_6 or k29_needs_bram_6 or k28_needs_bram_6 or k27_needs_bram_6 or k26_needs_bram_6 or k25_needs_bram_6 or k24_needs_bram_6) or ((k15_needs_bram_6 or k14_needs_bram_6 or k13_needs_bram_6 or k12_needs_bram_6 or k11_needs_bram_6 or k10_needs_bram_6 or k9_needs_bram_6 or k8_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6) and (not k18_needs_bram_6) and (not k19_needs_bram_6) and (not k20_needs_bram_6) and (not k21_needs_bram_6) and (not k22_needs_bram_6) and (not k23_needs_bram_6));
	bram_15_input_sel(3) <= (k31_needs_bram_7 or k30_needs_bram_7 or k29_needs_bram_7 or k28_needs_bram_7 or k27_needs_bram_7 or k26_needs_bram_7 or k25_needs_bram_7 or k24_needs_bram_7) or ((k15_needs_bram_7 or k14_needs_bram_7 or k13_needs_bram_7 or k12_needs_bram_7 or k11_needs_bram_7 or k10_needs_bram_7 or k9_needs_bram_7 or k8_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7) and (not k18_needs_bram_7) and (not k19_needs_bram_7) and (not k20_needs_bram_7) and (not k21_needs_bram_7) and (not k22_needs_bram_7) and (not k23_needs_bram_7));
	bram_17_input_sel(3) <= (k31_needs_bram_8 or k30_needs_bram_8 or k29_needs_bram_8 or k28_needs_bram_8 or k27_needs_bram_8 or k26_needs_bram_8 or k25_needs_bram_8 or k24_needs_bram_8) or ((k15_needs_bram_8 or k14_needs_bram_8 or k13_needs_bram_8 or k12_needs_bram_8 or k11_needs_bram_8 or k10_needs_bram_8 or k9_needs_bram_8 or k8_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8) and (not k18_needs_bram_8) and (not k19_needs_bram_8) and (not k20_needs_bram_8) and (not k21_needs_bram_8) and (not k22_needs_bram_8) and (not k23_needs_bram_8));
	bram_19_input_sel(3) <= (k31_needs_bram_9 or k30_needs_bram_9 or k29_needs_bram_9 or k28_needs_bram_9 or k27_needs_bram_9 or k26_needs_bram_9 or k25_needs_bram_9 or k24_needs_bram_9) or ((k15_needs_bram_9 or k14_needs_bram_9 or k13_needs_bram_9 or k12_needs_bram_9 or k11_needs_bram_9 or k10_needs_bram_9 or k9_needs_bram_9 or k8_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9) and (not k18_needs_bram_9) and (not k19_needs_bram_9) and (not k20_needs_bram_9) and (not k21_needs_bram_9) and (not k22_needs_bram_9) and (not k23_needs_bram_9));
	bram_21_input_sel(3) <= (k31_needs_bram_10 or k30_needs_bram_10 or k29_needs_bram_10 or k28_needs_bram_10 or k27_needs_bram_10 or k26_needs_bram_10 or k25_needs_bram_10 or k24_needs_bram_10) or ((k15_needs_bram_10 or k14_needs_bram_10 or k13_needs_bram_10 or k12_needs_bram_10 or k11_needs_bram_10 or k10_needs_bram_10 or k9_needs_bram_10 or k8_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10) and (not k18_needs_bram_10) and (not k19_needs_bram_10) and (not k20_needs_bram_10) and (not k21_needs_bram_10) and (not k22_needs_bram_10) and (not k23_needs_bram_10));
	bram_23_input_sel(3) <= (k31_needs_bram_11 or k30_needs_bram_11 or k29_needs_bram_11 or k28_needs_bram_11 or k27_needs_bram_11 or k26_needs_bram_11 or k25_needs_bram_11 or k24_needs_bram_11) or ((k15_needs_bram_11 or k14_needs_bram_11 or k13_needs_bram_11 or k12_needs_bram_11 or k11_needs_bram_11 or k10_needs_bram_11 or k9_needs_bram_11 or k8_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11) and (not k18_needs_bram_11) and (not k19_needs_bram_11) and (not k20_needs_bram_11) and (not k21_needs_bram_11) and (not k22_needs_bram_11) and (not k23_needs_bram_11));
	bram_25_input_sel(3) <= (k31_needs_bram_12 or k30_needs_bram_12 or k29_needs_bram_12 or k28_needs_bram_12 or k27_needs_bram_12 or k26_needs_bram_12 or k25_needs_bram_12 or k24_needs_bram_12) or ((k15_needs_bram_12 or k14_needs_bram_12 or k13_needs_bram_12 or k12_needs_bram_12 or k11_needs_bram_12 or k10_needs_bram_12 or k9_needs_bram_12 or k8_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12) and (not k18_needs_bram_12) and (not k19_needs_bram_12) and (not k20_needs_bram_12) and (not k21_needs_bram_12) and (not k22_needs_bram_12) and (not k23_needs_bram_12));
	bram_27_input_sel(3) <= (k31_needs_bram_13 or k30_needs_bram_13 or k29_needs_bram_13 or k28_needs_bram_13 or k27_needs_bram_13 or k26_needs_bram_13 or k25_needs_bram_13 or k24_needs_bram_13) or ((k15_needs_bram_13 or k14_needs_bram_13 or k13_needs_bram_13 or k12_needs_bram_13 or k11_needs_bram_13 or k10_needs_bram_13 or k9_needs_bram_13 or k8_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13) and (not k18_needs_bram_13) and (not k19_needs_bram_13) and (not k20_needs_bram_13) and (not k21_needs_bram_13) and (not k22_needs_bram_13) and (not k23_needs_bram_13));
	bram_29_input_sel(3) <= (k31_needs_bram_14 or k30_needs_bram_14 or k29_needs_bram_14 or k28_needs_bram_14 or k27_needs_bram_14 or k26_needs_bram_14 or k25_needs_bram_14 or k24_needs_bram_14) or ((k15_needs_bram_14 or k14_needs_bram_14 or k13_needs_bram_14 or k12_needs_bram_14 or k11_needs_bram_14 or k10_needs_bram_14 or k9_needs_bram_14 or k8_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14) and (not k18_needs_bram_14) and (not k19_needs_bram_14) and (not k20_needs_bram_14) and (not k21_needs_bram_14) and (not k22_needs_bram_14) and (not k23_needs_bram_14));
	bram_31_input_sel(3) <= (k31_needs_bram_15 or k30_needs_bram_15 or k29_needs_bram_15 or k28_needs_bram_15 or k27_needs_bram_15 or k26_needs_bram_15 or k25_needs_bram_15 or k24_needs_bram_15) or ((k15_needs_bram_15 or k14_needs_bram_15 or k13_needs_bram_15 or k12_needs_bram_15 or k11_needs_bram_15 or k10_needs_bram_15 or k9_needs_bram_15 or k8_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15) and (not k18_needs_bram_15) and (not k19_needs_bram_15) and (not k20_needs_bram_15) and (not k21_needs_bram_15) and (not k22_needs_bram_15) and (not k23_needs_bram_15));

	bram_1_input_sel(2) <= (k31_needs_bram_0 or k30_needs_bram_0 or k29_needs_bram_0 or k28_needs_bram_0) or ((k23_needs_bram_0 or k22_needs_bram_0 or k21_needs_bram_0 or k20_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k26_needs_bram_0) and (not k27_needs_bram_0)) or ((k15_needs_bram_0 or k14_needs_bram_0 or k13_needs_bram_0 or k12_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k26_needs_bram_0) and (not k27_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0) and (not k18_needs_bram_0) and (not k19_needs_bram_0)) or ((k7_needs_bram_0 or k6_needs_bram_0 or k5_needs_bram_0 or k4_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k26_needs_bram_0) and (not k27_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0) and (not k18_needs_bram_0) and (not k19_needs_bram_0) and (not k8_needs_bram_0) and (not k9_needs_bram_0) and (not k10_needs_bram_0) and (not k11_needs_bram_0));
	bram_3_input_sel(2) <= (k31_needs_bram_1 or k30_needs_bram_1 or k29_needs_bram_1 or k28_needs_bram_1) or ((k23_needs_bram_1 or k22_needs_bram_1 or k21_needs_bram_1 or k20_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k26_needs_bram_1) and (not k27_needs_bram_1)) or ((k15_needs_bram_1 or k14_needs_bram_1 or k13_needs_bram_1 or k12_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k26_needs_bram_1) and (not k27_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1) and (not k18_needs_bram_1) and (not k19_needs_bram_1)) or ((k7_needs_bram_1 or k6_needs_bram_1 or k5_needs_bram_1 or k4_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k26_needs_bram_1) and (not k27_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1) and (not k18_needs_bram_1) and (not k19_needs_bram_1) and (not k8_needs_bram_1) and (not k9_needs_bram_1) and (not k10_needs_bram_1) and (not k11_needs_bram_1));
	bram_5_input_sel(2) <= (k31_needs_bram_2 or k30_needs_bram_2 or k29_needs_bram_2 or k28_needs_bram_2) or ((k23_needs_bram_2 or k22_needs_bram_2 or k21_needs_bram_2 or k20_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k26_needs_bram_2) and (not k27_needs_bram_2)) or ((k15_needs_bram_2 or k14_needs_bram_2 or k13_needs_bram_2 or k12_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k26_needs_bram_2) and (not k27_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2) and (not k18_needs_bram_2) and (not k19_needs_bram_2)) or ((k7_needs_bram_2 or k6_needs_bram_2 or k5_needs_bram_2 or k4_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k26_needs_bram_2) and (not k27_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2) and (not k18_needs_bram_2) and (not k19_needs_bram_2) and (not k8_needs_bram_2) and (not k9_needs_bram_2) and (not k10_needs_bram_2) and (not k11_needs_bram_2));
	bram_7_input_sel(2) <= (k31_needs_bram_3 or k30_needs_bram_3 or k29_needs_bram_3 or k28_needs_bram_3) or ((k23_needs_bram_3 or k22_needs_bram_3 or k21_needs_bram_3 or k20_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k26_needs_bram_3) and (not k27_needs_bram_3)) or ((k15_needs_bram_3 or k14_needs_bram_3 or k13_needs_bram_3 or k12_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k26_needs_bram_3) and (not k27_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3) and (not k18_needs_bram_3) and (not k19_needs_bram_3)) or ((k7_needs_bram_3 or k6_needs_bram_3 or k5_needs_bram_3 or k4_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k26_needs_bram_3) and (not k27_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3) and (not k18_needs_bram_3) and (not k19_needs_bram_3) and (not k8_needs_bram_3) and (not k9_needs_bram_3) and (not k10_needs_bram_3) and (not k11_needs_bram_3));
	bram_9_input_sel(2) <= (k31_needs_bram_4 or k30_needs_bram_4 or k29_needs_bram_4 or k28_needs_bram_4) or ((k23_needs_bram_4 or k22_needs_bram_4 or k21_needs_bram_4 or k20_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k26_needs_bram_4) and (not k27_needs_bram_4)) or ((k15_needs_bram_4 or k14_needs_bram_4 or k13_needs_bram_4 or k12_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k26_needs_bram_4) and (not k27_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4) and (not k18_needs_bram_4) and (not k19_needs_bram_4)) or ((k7_needs_bram_4 or k6_needs_bram_4 or k5_needs_bram_4 or k4_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k26_needs_bram_4) and (not k27_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4) and (not k18_needs_bram_4) and (not k19_needs_bram_4) and (not k8_needs_bram_4) and (not k9_needs_bram_4) and (not k10_needs_bram_4) and (not k11_needs_bram_4));
	bram_11_input_sel(2) <= (k31_needs_bram_5 or k30_needs_bram_5 or k29_needs_bram_5 or k28_needs_bram_5) or ((k23_needs_bram_5 or k22_needs_bram_5 or k21_needs_bram_5 or k20_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k26_needs_bram_5) and (not k27_needs_bram_5)) or ((k15_needs_bram_5 or k14_needs_bram_5 or k13_needs_bram_5 or k12_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k26_needs_bram_5) and (not k27_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5) and (not k18_needs_bram_5) and (not k19_needs_bram_5)) or ((k7_needs_bram_5 or k6_needs_bram_5 or k5_needs_bram_5 or k4_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k26_needs_bram_5) and (not k27_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5) and (not k18_needs_bram_5) and (not k19_needs_bram_5) and (not k8_needs_bram_5) and (not k9_needs_bram_5) and (not k10_needs_bram_5) and (not k11_needs_bram_5));
	bram_13_input_sel(2) <= (k31_needs_bram_6 or k30_needs_bram_6 or k29_needs_bram_6 or k28_needs_bram_6) or ((k23_needs_bram_6 or k22_needs_bram_6 or k21_needs_bram_6 or k20_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k26_needs_bram_6) and (not k27_needs_bram_6)) or ((k15_needs_bram_6 or k14_needs_bram_6 or k13_needs_bram_6 or k12_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k26_needs_bram_6) and (not k27_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6) and (not k18_needs_bram_6) and (not k19_needs_bram_6)) or ((k7_needs_bram_6 or k6_needs_bram_6 or k5_needs_bram_6 or k4_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k26_needs_bram_6) and (not k27_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6) and (not k18_needs_bram_6) and (not k19_needs_bram_6) and (not k8_needs_bram_6) and (not k9_needs_bram_6) and (not k10_needs_bram_6) and (not k11_needs_bram_6));
	bram_15_input_sel(2) <= (k31_needs_bram_7 or k30_needs_bram_7 or k29_needs_bram_7 or k28_needs_bram_7) or ((k23_needs_bram_7 or k22_needs_bram_7 or k21_needs_bram_7 or k20_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k26_needs_bram_7) and (not k27_needs_bram_7)) or ((k15_needs_bram_7 or k14_needs_bram_7 or k13_needs_bram_7 or k12_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k26_needs_bram_7) and (not k27_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7) and (not k18_needs_bram_7) and (not k19_needs_bram_7)) or ((k7_needs_bram_7 or k6_needs_bram_7 or k5_needs_bram_7 or k4_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k26_needs_bram_7) and (not k27_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7) and (not k18_needs_bram_7) and (not k19_needs_bram_7) and (not k8_needs_bram_7) and (not k9_needs_bram_7) and (not k10_needs_bram_7) and (not k11_needs_bram_7));
	bram_17_input_sel(2) <= (k31_needs_bram_8 or k30_needs_bram_8 or k29_needs_bram_8 or k28_needs_bram_8) or ((k23_needs_bram_8 or k22_needs_bram_8 or k21_needs_bram_8 or k20_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k26_needs_bram_8) and (not k27_needs_bram_8)) or ((k15_needs_bram_8 or k14_needs_bram_8 or k13_needs_bram_8 or k12_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k26_needs_bram_8) and (not k27_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8) and (not k18_needs_bram_8) and (not k19_needs_bram_8)) or ((k7_needs_bram_8 or k6_needs_bram_8 or k5_needs_bram_8 or k4_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k26_needs_bram_8) and (not k27_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8) and (not k18_needs_bram_8) and (not k19_needs_bram_8) and (not k8_needs_bram_8) and (not k9_needs_bram_8) and (not k10_needs_bram_8) and (not k11_needs_bram_8));
	bram_19_input_sel(2) <= (k31_needs_bram_9 or k30_needs_bram_9 or k29_needs_bram_9 or k28_needs_bram_9) or ((k23_needs_bram_9 or k22_needs_bram_9 or k21_needs_bram_9 or k20_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k26_needs_bram_9) and (not k27_needs_bram_9)) or ((k15_needs_bram_9 or k14_needs_bram_9 or k13_needs_bram_9 or k12_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k26_needs_bram_9) and (not k27_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9) and (not k18_needs_bram_9) and (not k19_needs_bram_9)) or ((k7_needs_bram_9 or k6_needs_bram_9 or k5_needs_bram_9 or k4_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k26_needs_bram_9) and (not k27_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9) and (not k18_needs_bram_9) and (not k19_needs_bram_9) and (not k8_needs_bram_9) and (not k9_needs_bram_9) and (not k10_needs_bram_9) and (not k11_needs_bram_9));
	bram_21_input_sel(2) <= (k31_needs_bram_10 or k30_needs_bram_10 or k29_needs_bram_10 or k28_needs_bram_10) or ((k23_needs_bram_10 or k22_needs_bram_10 or k21_needs_bram_10 or k20_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k26_needs_bram_10) and (not k27_needs_bram_10)) or ((k15_needs_bram_10 or k14_needs_bram_10 or k13_needs_bram_10 or k12_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k26_needs_bram_10) and (not k27_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10) and (not k18_needs_bram_10) and (not k19_needs_bram_10)) or ((k7_needs_bram_10 or k6_needs_bram_10 or k5_needs_bram_10 or k4_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k26_needs_bram_10) and (not k27_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10) and (not k18_needs_bram_10) and (not k19_needs_bram_10) and (not k8_needs_bram_10) and (not k9_needs_bram_10) and (not k10_needs_bram_10) and (not k11_needs_bram_10));
	bram_23_input_sel(2) <= (k31_needs_bram_11 or k30_needs_bram_11 or k29_needs_bram_11 or k28_needs_bram_11) or ((k23_needs_bram_11 or k22_needs_bram_11 or k21_needs_bram_11 or k20_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k26_needs_bram_11) and (not k27_needs_bram_11)) or ((k15_needs_bram_11 or k14_needs_bram_11 or k13_needs_bram_11 or k12_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k26_needs_bram_11) and (not k27_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11) and (not k18_needs_bram_11) and (not k19_needs_bram_11)) or ((k7_needs_bram_11 or k6_needs_bram_11 or k5_needs_bram_11 or k4_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k26_needs_bram_11) and (not k27_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11) and (not k18_needs_bram_11) and (not k19_needs_bram_11) and (not k8_needs_bram_11) and (not k9_needs_bram_11) and (not k10_needs_bram_11) and (not k11_needs_bram_11));
	bram_25_input_sel(2) <= (k31_needs_bram_12 or k30_needs_bram_12 or k29_needs_bram_12 or k28_needs_bram_12) or ((k23_needs_bram_12 or k22_needs_bram_12 or k21_needs_bram_12 or k20_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k26_needs_bram_12) and (not k27_needs_bram_12)) or ((k15_needs_bram_12 or k14_needs_bram_12 or k13_needs_bram_12 or k12_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k26_needs_bram_12) and (not k27_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12) and (not k18_needs_bram_12) and (not k19_needs_bram_12)) or ((k7_needs_bram_12 or k6_needs_bram_12 or k5_needs_bram_12 or k4_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k26_needs_bram_12) and (not k27_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12) and (not k18_needs_bram_12) and (not k19_needs_bram_12) and (not k8_needs_bram_12) and (not k9_needs_bram_12) and (not k10_needs_bram_12) and (not k11_needs_bram_12));
	bram_27_input_sel(2) <= (k31_needs_bram_13 or k30_needs_bram_13 or k29_needs_bram_13 or k28_needs_bram_13) or ((k23_needs_bram_13 or k22_needs_bram_13 or k21_needs_bram_13 or k20_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k26_needs_bram_13) and (not k27_needs_bram_13)) or ((k15_needs_bram_13 or k14_needs_bram_13 or k13_needs_bram_13 or k12_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k26_needs_bram_13) and (not k27_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13) and (not k18_needs_bram_13) and (not k19_needs_bram_13)) or ((k7_needs_bram_13 or k6_needs_bram_13 or k5_needs_bram_13 or k4_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k26_needs_bram_13) and (not k27_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13) and (not k18_needs_bram_13) and (not k19_needs_bram_13) and (not k8_needs_bram_13) and (not k9_needs_bram_13) and (not k10_needs_bram_13) and (not k11_needs_bram_13));
	bram_29_input_sel(2) <= (k31_needs_bram_14 or k30_needs_bram_14 or k29_needs_bram_14 or k28_needs_bram_14) or ((k23_needs_bram_14 or k22_needs_bram_14 or k21_needs_bram_14 or k20_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k26_needs_bram_14) and (not k27_needs_bram_14)) or ((k15_needs_bram_14 or k14_needs_bram_14 or k13_needs_bram_14 or k12_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k26_needs_bram_14) and (not k27_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14) and (not k18_needs_bram_14) and (not k19_needs_bram_14)) or ((k7_needs_bram_14 or k6_needs_bram_14 or k5_needs_bram_14 or k4_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k26_needs_bram_14) and (not k27_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14) and (not k18_needs_bram_14) and (not k19_needs_bram_14) and (not k8_needs_bram_14) and (not k9_needs_bram_14) and (not k10_needs_bram_14) and (not k11_needs_bram_14));
	bram_31_input_sel(2) <= (k31_needs_bram_15 or k30_needs_bram_15 or k29_needs_bram_15 or k28_needs_bram_15) or ((k23_needs_bram_15 or k22_needs_bram_15 or k21_needs_bram_15 or k20_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k26_needs_bram_15) and (not k27_needs_bram_15)) or ((k15_needs_bram_15 or k14_needs_bram_15 or k13_needs_bram_15 or k12_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k26_needs_bram_15) and (not k27_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15) and (not k18_needs_bram_15) and (not k19_needs_bram_15)) or ((k7_needs_bram_15 or k6_needs_bram_15 or k5_needs_bram_15 or k4_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k26_needs_bram_15) and (not k27_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15) and (not k18_needs_bram_15) and (not k19_needs_bram_15) and (not k8_needs_bram_15) and (not k9_needs_bram_15) and (not k10_needs_bram_15) and (not k11_needs_bram_15));

	bram_1_input_sel(1) <= (k31_needs_bram_0 or k30_needs_bram_0) or ((k27_needs_bram_0 or k26_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0)) or ((k23_needs_bram_0 or k22_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0)) or ((k19_needs_bram_0 or k18_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k20_needs_bram_0) and (not k21_needs_bram_0)) or ((k15_needs_bram_0 or k14_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k20_needs_bram_0) and (not k21_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0)) or ((k11_needs_bram_0 or k10_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k20_needs_bram_0) and (not k21_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0) and (not k12_needs_bram_0) and (not k13_needs_bram_0)) or ((k7_needs_bram_0 or k6_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k20_needs_bram_0) and (not k21_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0) and (not k12_needs_bram_0) and (not k13_needs_bram_0) and (not k8_needs_bram_0) and (not k9_needs_bram_0)) or ((k3_needs_bram_0 or k2_needs_bram_0) and (not k28_needs_bram_0) and (not k29_needs_bram_0) and (not k24_needs_bram_0) and (not k25_needs_bram_0) and (not k20_needs_bram_0) and (not k21_needs_bram_0) and (not k16_needs_bram_0) and (not k17_needs_bram_0) and (not k12_needs_bram_0) and (not k13_needs_bram_0) and (not k8_needs_bram_0) and (not k9_needs_bram_0) and (not k4_needs_bram_0) and (not k5_needs_bram_0));
	bram_3_input_sel(1) <= (k31_needs_bram_1 or k30_needs_bram_1) or ((k27_needs_bram_1 or k26_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1)) or ((k23_needs_bram_1 or k22_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1)) or ((k19_needs_bram_1 or k18_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k20_needs_bram_1) and (not k21_needs_bram_1)) or ((k15_needs_bram_1 or k14_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k20_needs_bram_1) and (not k21_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1)) or ((k11_needs_bram_1 or k10_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k20_needs_bram_1) and (not k21_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1) and (not k12_needs_bram_1) and (not k13_needs_bram_1)) or ((k7_needs_bram_1 or k6_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k20_needs_bram_1) and (not k21_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1) and (not k12_needs_bram_1) and (not k13_needs_bram_1) and (not k8_needs_bram_1) and (not k9_needs_bram_1)) or ((k3_needs_bram_1 or k2_needs_bram_1) and (not k28_needs_bram_1) and (not k29_needs_bram_1) and (not k24_needs_bram_1) and (not k25_needs_bram_1) and (not k20_needs_bram_1) and (not k21_needs_bram_1) and (not k16_needs_bram_1) and (not k17_needs_bram_1) and (not k12_needs_bram_1) and (not k13_needs_bram_1) and (not k8_needs_bram_1) and (not k9_needs_bram_1) and (not k4_needs_bram_1) and (not k5_needs_bram_1));
	bram_5_input_sel(1) <= (k31_needs_bram_2 or k30_needs_bram_2) or ((k27_needs_bram_2 or k26_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2)) or ((k23_needs_bram_2 or k22_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2)) or ((k19_needs_bram_2 or k18_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k20_needs_bram_2) and (not k21_needs_bram_2)) or ((k15_needs_bram_2 or k14_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k20_needs_bram_2) and (not k21_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2)) or ((k11_needs_bram_2 or k10_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k20_needs_bram_2) and (not k21_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2) and (not k12_needs_bram_2) and (not k13_needs_bram_2)) or ((k7_needs_bram_2 or k6_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k20_needs_bram_2) and (not k21_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2) and (not k12_needs_bram_2) and (not k13_needs_bram_2) and (not k8_needs_bram_2) and (not k9_needs_bram_2)) or ((k3_needs_bram_2 or k2_needs_bram_2) and (not k28_needs_bram_2) and (not k29_needs_bram_2) and (not k24_needs_bram_2) and (not k25_needs_bram_2) and (not k20_needs_bram_2) and (not k21_needs_bram_2) and (not k16_needs_bram_2) and (not k17_needs_bram_2) and (not k12_needs_bram_2) and (not k13_needs_bram_2) and (not k8_needs_bram_2) and (not k9_needs_bram_2) and (not k4_needs_bram_2) and (not k5_needs_bram_2));
	bram_7_input_sel(1) <= (k31_needs_bram_3 or k30_needs_bram_3) or ((k27_needs_bram_3 or k26_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3)) or ((k23_needs_bram_3 or k22_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3)) or ((k19_needs_bram_3 or k18_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k20_needs_bram_3) and (not k21_needs_bram_3)) or ((k15_needs_bram_3 or k14_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k20_needs_bram_3) and (not k21_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3)) or ((k11_needs_bram_3 or k10_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k20_needs_bram_3) and (not k21_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3) and (not k12_needs_bram_3) and (not k13_needs_bram_3)) or ((k7_needs_bram_3 or k6_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k20_needs_bram_3) and (not k21_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3) and (not k12_needs_bram_3) and (not k13_needs_bram_3) and (not k8_needs_bram_3) and (not k9_needs_bram_3)) or ((k3_needs_bram_3 or k2_needs_bram_3) and (not k28_needs_bram_3) and (not k29_needs_bram_3) and (not k24_needs_bram_3) and (not k25_needs_bram_3) and (not k20_needs_bram_3) and (not k21_needs_bram_3) and (not k16_needs_bram_3) and (not k17_needs_bram_3) and (not k12_needs_bram_3) and (not k13_needs_bram_3) and (not k8_needs_bram_3) and (not k9_needs_bram_3) and (not k4_needs_bram_3) and (not k5_needs_bram_3));
	bram_9_input_sel(1) <= (k31_needs_bram_4 or k30_needs_bram_4) or ((k27_needs_bram_4 or k26_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4)) or ((k23_needs_bram_4 or k22_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4)) or ((k19_needs_bram_4 or k18_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k20_needs_bram_4) and (not k21_needs_bram_4)) or ((k15_needs_bram_4 or k14_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k20_needs_bram_4) and (not k21_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4)) or ((k11_needs_bram_4 or k10_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k20_needs_bram_4) and (not k21_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4) and (not k12_needs_bram_4) and (not k13_needs_bram_4)) or ((k7_needs_bram_4 or k6_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k20_needs_bram_4) and (not k21_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4) and (not k12_needs_bram_4) and (not k13_needs_bram_4) and (not k8_needs_bram_4) and (not k9_needs_bram_4)) or ((k3_needs_bram_4 or k2_needs_bram_4) and (not k28_needs_bram_4) and (not k29_needs_bram_4) and (not k24_needs_bram_4) and (not k25_needs_bram_4) and (not k20_needs_bram_4) and (not k21_needs_bram_4) and (not k16_needs_bram_4) and (not k17_needs_bram_4) and (not k12_needs_bram_4) and (not k13_needs_bram_4) and (not k8_needs_bram_4) and (not k9_needs_bram_4) and (not k4_needs_bram_4) and (not k5_needs_bram_4));
	bram_11_input_sel(1) <= (k31_needs_bram_5 or k30_needs_bram_5) or ((k27_needs_bram_5 or k26_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5)) or ((k23_needs_bram_5 or k22_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5)) or ((k19_needs_bram_5 or k18_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k20_needs_bram_5) and (not k21_needs_bram_5)) or ((k15_needs_bram_5 or k14_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k20_needs_bram_5) and (not k21_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5)) or ((k11_needs_bram_5 or k10_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k20_needs_bram_5) and (not k21_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5) and (not k12_needs_bram_5) and (not k13_needs_bram_5)) or ((k7_needs_bram_5 or k6_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k20_needs_bram_5) and (not k21_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5) and (not k12_needs_bram_5) and (not k13_needs_bram_5) and (not k8_needs_bram_5) and (not k9_needs_bram_5)) or ((k3_needs_bram_5 or k2_needs_bram_5) and (not k28_needs_bram_5) and (not k29_needs_bram_5) and (not k24_needs_bram_5) and (not k25_needs_bram_5) and (not k20_needs_bram_5) and (not k21_needs_bram_5) and (not k16_needs_bram_5) and (not k17_needs_bram_5) and (not k12_needs_bram_5) and (not k13_needs_bram_5) and (not k8_needs_bram_5) and (not k9_needs_bram_5) and (not k4_needs_bram_5) and (not k5_needs_bram_5));
	bram_13_input_sel(1) <= (k31_needs_bram_6 or k30_needs_bram_6) or ((k27_needs_bram_6 or k26_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6)) or ((k23_needs_bram_6 or k22_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6)) or ((k19_needs_bram_6 or k18_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k20_needs_bram_6) and (not k21_needs_bram_6)) or ((k15_needs_bram_6 or k14_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k20_needs_bram_6) and (not k21_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6)) or ((k11_needs_bram_6 or k10_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k20_needs_bram_6) and (not k21_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6) and (not k12_needs_bram_6) and (not k13_needs_bram_6)) or ((k7_needs_bram_6 or k6_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k20_needs_bram_6) and (not k21_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6) and (not k12_needs_bram_6) and (not k13_needs_bram_6) and (not k8_needs_bram_6) and (not k9_needs_bram_6)) or ((k3_needs_bram_6 or k2_needs_bram_6) and (not k28_needs_bram_6) and (not k29_needs_bram_6) and (not k24_needs_bram_6) and (not k25_needs_bram_6) and (not k20_needs_bram_6) and (not k21_needs_bram_6) and (not k16_needs_bram_6) and (not k17_needs_bram_6) and (not k12_needs_bram_6) and (not k13_needs_bram_6) and (not k8_needs_bram_6) and (not k9_needs_bram_6) and (not k4_needs_bram_6) and (not k5_needs_bram_6));
	bram_15_input_sel(1) <= (k31_needs_bram_7 or k30_needs_bram_7) or ((k27_needs_bram_7 or k26_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7)) or ((k23_needs_bram_7 or k22_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7)) or ((k19_needs_bram_7 or k18_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k20_needs_bram_7) and (not k21_needs_bram_7)) or ((k15_needs_bram_7 or k14_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k20_needs_bram_7) and (not k21_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7)) or ((k11_needs_bram_7 or k10_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k20_needs_bram_7) and (not k21_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7) and (not k12_needs_bram_7) and (not k13_needs_bram_7)) or ((k7_needs_bram_7 or k6_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k20_needs_bram_7) and (not k21_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7) and (not k12_needs_bram_7) and (not k13_needs_bram_7) and (not k8_needs_bram_7) and (not k9_needs_bram_7)) or ((k3_needs_bram_7 or k2_needs_bram_7) and (not k28_needs_bram_7) and (not k29_needs_bram_7) and (not k24_needs_bram_7) and (not k25_needs_bram_7) and (not k20_needs_bram_7) and (not k21_needs_bram_7) and (not k16_needs_bram_7) and (not k17_needs_bram_7) and (not k12_needs_bram_7) and (not k13_needs_bram_7) and (not k8_needs_bram_7) and (not k9_needs_bram_7) and (not k4_needs_bram_7) and (not k5_needs_bram_7));
	bram_17_input_sel(1) <= (k31_needs_bram_8 or k30_needs_bram_8) or ((k27_needs_bram_8 or k26_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8)) or ((k23_needs_bram_8 or k22_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8)) or ((k19_needs_bram_8 or k18_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k20_needs_bram_8) and (not k21_needs_bram_8)) or ((k15_needs_bram_8 or k14_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k20_needs_bram_8) and (not k21_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8)) or ((k11_needs_bram_8 or k10_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k20_needs_bram_8) and (not k21_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8) and (not k12_needs_bram_8) and (not k13_needs_bram_8)) or ((k7_needs_bram_8 or k6_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k20_needs_bram_8) and (not k21_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8) and (not k12_needs_bram_8) and (not k13_needs_bram_8) and (not k8_needs_bram_8) and (not k9_needs_bram_8)) or ((k3_needs_bram_8 or k2_needs_bram_8) and (not k28_needs_bram_8) and (not k29_needs_bram_8) and (not k24_needs_bram_8) and (not k25_needs_bram_8) and (not k20_needs_bram_8) and (not k21_needs_bram_8) and (not k16_needs_bram_8) and (not k17_needs_bram_8) and (not k12_needs_bram_8) and (not k13_needs_bram_8) and (not k8_needs_bram_8) and (not k9_needs_bram_8) and (not k4_needs_bram_8) and (not k5_needs_bram_8));
	bram_19_input_sel(1) <= (k31_needs_bram_9 or k30_needs_bram_9) or ((k27_needs_bram_9 or k26_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9)) or ((k23_needs_bram_9 or k22_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9)) or ((k19_needs_bram_9 or k18_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k20_needs_bram_9) and (not k21_needs_bram_9)) or ((k15_needs_bram_9 or k14_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k20_needs_bram_9) and (not k21_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9)) or ((k11_needs_bram_9 or k10_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k20_needs_bram_9) and (not k21_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9) and (not k12_needs_bram_9) and (not k13_needs_bram_9)) or ((k7_needs_bram_9 or k6_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k20_needs_bram_9) and (not k21_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9) and (not k12_needs_bram_9) and (not k13_needs_bram_9) and (not k8_needs_bram_9) and (not k9_needs_bram_9)) or ((k3_needs_bram_9 or k2_needs_bram_9) and (not k28_needs_bram_9) and (not k29_needs_bram_9) and (not k24_needs_bram_9) and (not k25_needs_bram_9) and (not k20_needs_bram_9) and (not k21_needs_bram_9) and (not k16_needs_bram_9) and (not k17_needs_bram_9) and (not k12_needs_bram_9) and (not k13_needs_bram_9) and (not k8_needs_bram_9) and (not k9_needs_bram_9) and (not k4_needs_bram_9) and (not k5_needs_bram_9));
	bram_21_input_sel(1) <= (k31_needs_bram_10 or k30_needs_bram_10) or ((k27_needs_bram_10 or k26_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10)) or ((k23_needs_bram_10 or k22_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10)) or ((k19_needs_bram_10 or k18_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k20_needs_bram_10) and (not k21_needs_bram_10)) or ((k15_needs_bram_10 or k14_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k20_needs_bram_10) and (not k21_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10)) or ((k11_needs_bram_10 or k10_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k20_needs_bram_10) and (not k21_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10) and (not k12_needs_bram_10) and (not k13_needs_bram_10)) or ((k7_needs_bram_10 or k6_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k20_needs_bram_10) and (not k21_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10) and (not k12_needs_bram_10) and (not k13_needs_bram_10) and (not k8_needs_bram_10) and (not k9_needs_bram_10)) or ((k3_needs_bram_10 or k2_needs_bram_10) and (not k28_needs_bram_10) and (not k29_needs_bram_10) and (not k24_needs_bram_10) and (not k25_needs_bram_10) and (not k20_needs_bram_10) and (not k21_needs_bram_10) and (not k16_needs_bram_10) and (not k17_needs_bram_10) and (not k12_needs_bram_10) and (not k13_needs_bram_10) and (not k8_needs_bram_10) and (not k9_needs_bram_10) and (not k4_needs_bram_10) and (not k5_needs_bram_10));
	bram_23_input_sel(1) <= (k31_needs_bram_11 or k30_needs_bram_11) or ((k27_needs_bram_11 or k26_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11)) or ((k23_needs_bram_11 or k22_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11)) or ((k19_needs_bram_11 or k18_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k20_needs_bram_11) and (not k21_needs_bram_11)) or ((k15_needs_bram_11 or k14_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k20_needs_bram_11) and (not k21_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11)) or ((k11_needs_bram_11 or k10_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k20_needs_bram_11) and (not k21_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11) and (not k12_needs_bram_11) and (not k13_needs_bram_11)) or ((k7_needs_bram_11 or k6_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k20_needs_bram_11) and (not k21_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11) and (not k12_needs_bram_11) and (not k13_needs_bram_11) and (not k8_needs_bram_11) and (not k9_needs_bram_11)) or ((k3_needs_bram_11 or k2_needs_bram_11) and (not k28_needs_bram_11) and (not k29_needs_bram_11) and (not k24_needs_bram_11) and (not k25_needs_bram_11) and (not k20_needs_bram_11) and (not k21_needs_bram_11) and (not k16_needs_bram_11) and (not k17_needs_bram_11) and (not k12_needs_bram_11) and (not k13_needs_bram_11) and (not k8_needs_bram_11) and (not k9_needs_bram_11) and (not k4_needs_bram_11) and (not k5_needs_bram_11));
	bram_25_input_sel(1) <= (k31_needs_bram_12 or k30_needs_bram_12) or ((k27_needs_bram_12 or k26_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12)) or ((k23_needs_bram_12 or k22_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12)) or ((k19_needs_bram_12 or k18_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k20_needs_bram_12) and (not k21_needs_bram_12)) or ((k15_needs_bram_12 or k14_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k20_needs_bram_12) and (not k21_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12)) or ((k11_needs_bram_12 or k10_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k20_needs_bram_12) and (not k21_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12) and (not k12_needs_bram_12) and (not k13_needs_bram_12)) or ((k7_needs_bram_12 or k6_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k20_needs_bram_12) and (not k21_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12) and (not k12_needs_bram_12) and (not k13_needs_bram_12) and (not k8_needs_bram_12) and (not k9_needs_bram_12)) or ((k3_needs_bram_12 or k2_needs_bram_12) and (not k28_needs_bram_12) and (not k29_needs_bram_12) and (not k24_needs_bram_12) and (not k25_needs_bram_12) and (not k20_needs_bram_12) and (not k21_needs_bram_12) and (not k16_needs_bram_12) and (not k17_needs_bram_12) and (not k12_needs_bram_12) and (not k13_needs_bram_12) and (not k8_needs_bram_12) and (not k9_needs_bram_12) and (not k4_needs_bram_12) and (not k5_needs_bram_12));
	bram_27_input_sel(1) <= (k31_needs_bram_13 or k30_needs_bram_13) or ((k27_needs_bram_13 or k26_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13)) or ((k23_needs_bram_13 or k22_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13)) or ((k19_needs_bram_13 or k18_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k20_needs_bram_13) and (not k21_needs_bram_13)) or ((k15_needs_bram_13 or k14_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k20_needs_bram_13) and (not k21_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13)) or ((k11_needs_bram_13 or k10_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k20_needs_bram_13) and (not k21_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13) and (not k12_needs_bram_13) and (not k13_needs_bram_13)) or ((k7_needs_bram_13 or k6_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k20_needs_bram_13) and (not k21_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13) and (not k12_needs_bram_13) and (not k13_needs_bram_13) and (not k8_needs_bram_13) and (not k9_needs_bram_13)) or ((k3_needs_bram_13 or k2_needs_bram_13) and (not k28_needs_bram_13) and (not k29_needs_bram_13) and (not k24_needs_bram_13) and (not k25_needs_bram_13) and (not k20_needs_bram_13) and (not k21_needs_bram_13) and (not k16_needs_bram_13) and (not k17_needs_bram_13) and (not k12_needs_bram_13) and (not k13_needs_bram_13) and (not k8_needs_bram_13) and (not k9_needs_bram_13) and (not k4_needs_bram_13) and (not k5_needs_bram_13));
	bram_29_input_sel(1) <= (k31_needs_bram_14 or k30_needs_bram_14) or ((k27_needs_bram_14 or k26_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14)) or ((k23_needs_bram_14 or k22_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14)) or ((k19_needs_bram_14 or k18_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k20_needs_bram_14) and (not k21_needs_bram_14)) or ((k15_needs_bram_14 or k14_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k20_needs_bram_14) and (not k21_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14)) or ((k11_needs_bram_14 or k10_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k20_needs_bram_14) and (not k21_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14) and (not k12_needs_bram_14) and (not k13_needs_bram_14)) or ((k7_needs_bram_14 or k6_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k20_needs_bram_14) and (not k21_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14) and (not k12_needs_bram_14) and (not k13_needs_bram_14) and (not k8_needs_bram_14) and (not k9_needs_bram_14)) or ((k3_needs_bram_14 or k2_needs_bram_14) and (not k28_needs_bram_14) and (not k29_needs_bram_14) and (not k24_needs_bram_14) and (not k25_needs_bram_14) and (not k20_needs_bram_14) and (not k21_needs_bram_14) and (not k16_needs_bram_14) and (not k17_needs_bram_14) and (not k12_needs_bram_14) and (not k13_needs_bram_14) and (not k8_needs_bram_14) and (not k9_needs_bram_14) and (not k4_needs_bram_14) and (not k5_needs_bram_14));
	bram_31_input_sel(1) <= (k31_needs_bram_15 or k30_needs_bram_15) or ((k27_needs_bram_15 or k26_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15)) or ((k23_needs_bram_15 or k22_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15)) or ((k19_needs_bram_15 or k18_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k20_needs_bram_15) and (not k21_needs_bram_15)) or ((k15_needs_bram_15 or k14_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k20_needs_bram_15) and (not k21_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15)) or ((k11_needs_bram_15 or k10_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k20_needs_bram_15) and (not k21_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15) and (not k12_needs_bram_15) and (not k13_needs_bram_15)) or ((k7_needs_bram_15 or k6_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k20_needs_bram_15) and (not k21_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15) and (not k12_needs_bram_15) and (not k13_needs_bram_15) and (not k8_needs_bram_15) and (not k9_needs_bram_15)) or ((k3_needs_bram_15 or k2_needs_bram_15) and (not k28_needs_bram_15) and (not k29_needs_bram_15) and (not k24_needs_bram_15) and (not k25_needs_bram_15) and (not k20_needs_bram_15) and (not k21_needs_bram_15) and (not k16_needs_bram_15) and (not k17_needs_bram_15) and (not k12_needs_bram_15) and (not k13_needs_bram_15) and (not k8_needs_bram_15) and (not k9_needs_bram_15) and (not k4_needs_bram_15) and (not k5_needs_bram_15));

	bram_1_input_sel(0) <= (k31_needs_bram_0) or ((k29_needs_bram_0) and (not k30_needs_bram_0)) or ((k27_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0)) or ((k25_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0)) or ((k23_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0)) or ((k21_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0)) or ((k19_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0)) or ((k17_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0)) or ((k15_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0)) or ((k13_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0)) or ((k11_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0) and (not k12_needs_bram_0)) or ((k9_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0) and (not k12_needs_bram_0) and (not k10_needs_bram_0)) or ((k7_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0) and (not k12_needs_bram_0) and (not k10_needs_bram_0) and (not k8_needs_bram_0)) or ((k5_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0) and (not k12_needs_bram_0) and (not k10_needs_bram_0) and (not k8_needs_bram_0) and (not k6_needs_bram_0)) or ((k3_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0) and (not k12_needs_bram_0) and (not k10_needs_bram_0) and (not k8_needs_bram_0) and (not k6_needs_bram_0) and (not k4_needs_bram_0)) or ((k1_needs_bram_0) and (not k30_needs_bram_0) and (not k28_needs_bram_0) and (not k26_needs_bram_0) and (not k24_needs_bram_0) and (not k22_needs_bram_0) and (not k20_needs_bram_0) and (not k18_needs_bram_0) and (not k16_needs_bram_0) and (not k14_needs_bram_0) and (not k12_needs_bram_0) and (not k10_needs_bram_0) and (not k8_needs_bram_0) and (not k6_needs_bram_0) and (not k4_needs_bram_0) and (not k2_needs_bram_0));
	bram_3_input_sel(0) <= (k31_needs_bram_1) or ((k29_needs_bram_1) and (not k30_needs_bram_1)) or ((k27_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1)) or ((k25_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1)) or ((k23_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1)) or ((k21_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1)) or ((k19_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1)) or ((k17_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1)) or ((k15_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1)) or ((k13_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1)) or ((k11_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1) and (not k12_needs_bram_1)) or ((k9_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1) and (not k12_needs_bram_1) and (not k10_needs_bram_1)) or ((k7_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1) and (not k12_needs_bram_1) and (not k10_needs_bram_1) and (not k8_needs_bram_1)) or ((k5_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1) and (not k12_needs_bram_1) and (not k10_needs_bram_1) and (not k8_needs_bram_1) and (not k6_needs_bram_1)) or ((k3_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1) and (not k12_needs_bram_1) and (not k10_needs_bram_1) and (not k8_needs_bram_1) and (not k6_needs_bram_1) and (not k4_needs_bram_1)) or ((k1_needs_bram_1) and (not k30_needs_bram_1) and (not k28_needs_bram_1) and (not k26_needs_bram_1) and (not k24_needs_bram_1) and (not k22_needs_bram_1) and (not k20_needs_bram_1) and (not k18_needs_bram_1) and (not k16_needs_bram_1) and (not k14_needs_bram_1) and (not k12_needs_bram_1) and (not k10_needs_bram_1) and (not k8_needs_bram_1) and (not k6_needs_bram_1) and (not k4_needs_bram_1) and (not k2_needs_bram_1));
	bram_5_input_sel(0) <= (k31_needs_bram_2) or ((k29_needs_bram_2) and (not k30_needs_bram_2)) or ((k27_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2)) or ((k25_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2)) or ((k23_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2)) or ((k21_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2)) or ((k19_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2)) or ((k17_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2)) or ((k15_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2)) or ((k13_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2)) or ((k11_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2) and (not k12_needs_bram_2)) or ((k9_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2) and (not k12_needs_bram_2) and (not k10_needs_bram_2)) or ((k7_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2) and (not k12_needs_bram_2) and (not k10_needs_bram_2) and (not k8_needs_bram_2)) or ((k5_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2) and (not k12_needs_bram_2) and (not k10_needs_bram_2) and (not k8_needs_bram_2) and (not k6_needs_bram_2)) or ((k3_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2) and (not k12_needs_bram_2) and (not k10_needs_bram_2) and (not k8_needs_bram_2) and (not k6_needs_bram_2) and (not k4_needs_bram_2)) or ((k1_needs_bram_2) and (not k30_needs_bram_2) and (not k28_needs_bram_2) and (not k26_needs_bram_2) and (not k24_needs_bram_2) and (not k22_needs_bram_2) and (not k20_needs_bram_2) and (not k18_needs_bram_2) and (not k16_needs_bram_2) and (not k14_needs_bram_2) and (not k12_needs_bram_2) and (not k10_needs_bram_2) and (not k8_needs_bram_2) and (not k6_needs_bram_2) and (not k4_needs_bram_2) and (not k2_needs_bram_2));
	bram_7_input_sel(0) <= (k31_needs_bram_3) or ((k29_needs_bram_3) and (not k30_needs_bram_3)) or ((k27_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3)) or ((k25_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3)) or ((k23_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3)) or ((k21_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3)) or ((k19_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3)) or ((k17_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3)) or ((k15_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3)) or ((k13_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3)) or ((k11_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3) and (not k12_needs_bram_3)) or ((k9_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3) and (not k12_needs_bram_3) and (not k10_needs_bram_3)) or ((k7_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3) and (not k12_needs_bram_3) and (not k10_needs_bram_3) and (not k8_needs_bram_3)) or ((k5_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3) and (not k12_needs_bram_3) and (not k10_needs_bram_3) and (not k8_needs_bram_3) and (not k6_needs_bram_3)) or ((k3_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3) and (not k12_needs_bram_3) and (not k10_needs_bram_3) and (not k8_needs_bram_3) and (not k6_needs_bram_3) and (not k4_needs_bram_3)) or ((k1_needs_bram_3) and (not k30_needs_bram_3) and (not k28_needs_bram_3) and (not k26_needs_bram_3) and (not k24_needs_bram_3) and (not k22_needs_bram_3) and (not k20_needs_bram_3) and (not k18_needs_bram_3) and (not k16_needs_bram_3) and (not k14_needs_bram_3) and (not k12_needs_bram_3) and (not k10_needs_bram_3) and (not k8_needs_bram_3) and (not k6_needs_bram_3) and (not k4_needs_bram_3) and (not k2_needs_bram_3));
	bram_9_input_sel(0) <= (k31_needs_bram_4) or ((k29_needs_bram_4) and (not k30_needs_bram_4)) or ((k27_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4)) or ((k25_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4)) or ((k23_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4)) or ((k21_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4)) or ((k19_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4)) or ((k17_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4)) or ((k15_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4)) or ((k13_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4)) or ((k11_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4) and (not k12_needs_bram_4)) or ((k9_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4) and (not k12_needs_bram_4) and (not k10_needs_bram_4)) or ((k7_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4) and (not k12_needs_bram_4) and (not k10_needs_bram_4) and (not k8_needs_bram_4)) or ((k5_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4) and (not k12_needs_bram_4) and (not k10_needs_bram_4) and (not k8_needs_bram_4) and (not k6_needs_bram_4)) or ((k3_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4) and (not k12_needs_bram_4) and (not k10_needs_bram_4) and (not k8_needs_bram_4) and (not k6_needs_bram_4) and (not k4_needs_bram_4)) or ((k1_needs_bram_4) and (not k30_needs_bram_4) and (not k28_needs_bram_4) and (not k26_needs_bram_4) and (not k24_needs_bram_4) and (not k22_needs_bram_4) and (not k20_needs_bram_4) and (not k18_needs_bram_4) and (not k16_needs_bram_4) and (not k14_needs_bram_4) and (not k12_needs_bram_4) and (not k10_needs_bram_4) and (not k8_needs_bram_4) and (not k6_needs_bram_4) and (not k4_needs_bram_4) and (not k2_needs_bram_4));
	bram_11_input_sel(0) <= (k31_needs_bram_5) or ((k29_needs_bram_5) and (not k30_needs_bram_5)) or ((k27_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5)) or ((k25_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5)) or ((k23_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5)) or ((k21_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5)) or ((k19_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5)) or ((k17_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5)) or ((k15_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5)) or ((k13_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5)) or ((k11_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5) and (not k12_needs_bram_5)) or ((k9_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5) and (not k12_needs_bram_5) and (not k10_needs_bram_5)) or ((k7_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5) and (not k12_needs_bram_5) and (not k10_needs_bram_5) and (not k8_needs_bram_5)) or ((k5_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5) and (not k12_needs_bram_5) and (not k10_needs_bram_5) and (not k8_needs_bram_5) and (not k6_needs_bram_5)) or ((k3_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5) and (not k12_needs_bram_5) and (not k10_needs_bram_5) and (not k8_needs_bram_5) and (not k6_needs_bram_5) and (not k4_needs_bram_5)) or ((k1_needs_bram_5) and (not k30_needs_bram_5) and (not k28_needs_bram_5) and (not k26_needs_bram_5) and (not k24_needs_bram_5) and (not k22_needs_bram_5) and (not k20_needs_bram_5) and (not k18_needs_bram_5) and (not k16_needs_bram_5) and (not k14_needs_bram_5) and (not k12_needs_bram_5) and (not k10_needs_bram_5) and (not k8_needs_bram_5) and (not k6_needs_bram_5) and (not k4_needs_bram_5) and (not k2_needs_bram_5));
	bram_13_input_sel(0) <= (k31_needs_bram_6) or ((k29_needs_bram_6) and (not k30_needs_bram_6)) or ((k27_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6)) or ((k25_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6)) or ((k23_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6)) or ((k21_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6)) or ((k19_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6)) or ((k17_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6)) or ((k15_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6)) or ((k13_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6)) or ((k11_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6) and (not k12_needs_bram_6)) or ((k9_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6) and (not k12_needs_bram_6) and (not k10_needs_bram_6)) or ((k7_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6) and (not k12_needs_bram_6) and (not k10_needs_bram_6) and (not k8_needs_bram_6)) or ((k5_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6) and (not k12_needs_bram_6) and (not k10_needs_bram_6) and (not k8_needs_bram_6) and (not k6_needs_bram_6)) or ((k3_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6) and (not k12_needs_bram_6) and (not k10_needs_bram_6) and (not k8_needs_bram_6) and (not k6_needs_bram_6) and (not k4_needs_bram_6)) or ((k1_needs_bram_6) and (not k30_needs_bram_6) and (not k28_needs_bram_6) and (not k26_needs_bram_6) and (not k24_needs_bram_6) and (not k22_needs_bram_6) and (not k20_needs_bram_6) and (not k18_needs_bram_6) and (not k16_needs_bram_6) and (not k14_needs_bram_6) and (not k12_needs_bram_6) and (not k10_needs_bram_6) and (not k8_needs_bram_6) and (not k6_needs_bram_6) and (not k4_needs_bram_6) and (not k2_needs_bram_6));
	bram_15_input_sel(0) <= (k31_needs_bram_7) or ((k29_needs_bram_7) and (not k30_needs_bram_7)) or ((k27_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7)) or ((k25_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7)) or ((k23_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7)) or ((k21_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7)) or ((k19_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7)) or ((k17_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7)) or ((k15_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7)) or ((k13_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7)) or ((k11_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7) and (not k12_needs_bram_7)) or ((k9_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7) and (not k12_needs_bram_7) and (not k10_needs_bram_7)) or ((k7_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7) and (not k12_needs_bram_7) and (not k10_needs_bram_7) and (not k8_needs_bram_7)) or ((k5_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7) and (not k12_needs_bram_7) and (not k10_needs_bram_7) and (not k8_needs_bram_7) and (not k6_needs_bram_7)) or ((k3_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7) and (not k12_needs_bram_7) and (not k10_needs_bram_7) and (not k8_needs_bram_7) and (not k6_needs_bram_7) and (not k4_needs_bram_7)) or ((k1_needs_bram_7) and (not k30_needs_bram_7) and (not k28_needs_bram_7) and (not k26_needs_bram_7) and (not k24_needs_bram_7) and (not k22_needs_bram_7) and (not k20_needs_bram_7) and (not k18_needs_bram_7) and (not k16_needs_bram_7) and (not k14_needs_bram_7) and (not k12_needs_bram_7) and (not k10_needs_bram_7) and (not k8_needs_bram_7) and (not k6_needs_bram_7) and (not k4_needs_bram_7) and (not k2_needs_bram_7));
	bram_17_input_sel(0) <= (k31_needs_bram_8) or ((k29_needs_bram_8) and (not k30_needs_bram_8)) or ((k27_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8)) or ((k25_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8)) or ((k23_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8)) or ((k21_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8)) or ((k19_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8)) or ((k17_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8)) or ((k15_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8)) or ((k13_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8)) or ((k11_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8) and (not k12_needs_bram_8)) or ((k9_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8) and (not k12_needs_bram_8) and (not k10_needs_bram_8)) or ((k7_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8) and (not k12_needs_bram_8) and (not k10_needs_bram_8) and (not k8_needs_bram_8)) or ((k5_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8) and (not k12_needs_bram_8) and (not k10_needs_bram_8) and (not k8_needs_bram_8) and (not k6_needs_bram_8)) or ((k3_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8) and (not k12_needs_bram_8) and (not k10_needs_bram_8) and (not k8_needs_bram_8) and (not k6_needs_bram_8) and (not k4_needs_bram_8)) or ((k1_needs_bram_8) and (not k30_needs_bram_8) and (not k28_needs_bram_8) and (not k26_needs_bram_8) and (not k24_needs_bram_8) and (not k22_needs_bram_8) and (not k20_needs_bram_8) and (not k18_needs_bram_8) and (not k16_needs_bram_8) and (not k14_needs_bram_8) and (not k12_needs_bram_8) and (not k10_needs_bram_8) and (not k8_needs_bram_8) and (not k6_needs_bram_8) and (not k4_needs_bram_8) and (not k2_needs_bram_8));
	bram_19_input_sel(0) <= (k31_needs_bram_9) or ((k29_needs_bram_9) and (not k30_needs_bram_9)) or ((k27_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9)) or ((k25_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9)) or ((k23_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9)) or ((k21_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9)) or ((k19_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9)) or ((k17_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9)) or ((k15_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9)) or ((k13_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9)) or ((k11_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9) and (not k12_needs_bram_9)) or ((k9_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9) and (not k12_needs_bram_9) and (not k10_needs_bram_9)) or ((k7_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9) and (not k12_needs_bram_9) and (not k10_needs_bram_9) and (not k8_needs_bram_9)) or ((k5_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9) and (not k12_needs_bram_9) and (not k10_needs_bram_9) and (not k8_needs_bram_9) and (not k6_needs_bram_9)) or ((k3_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9) and (not k12_needs_bram_9) and (not k10_needs_bram_9) and (not k8_needs_bram_9) and (not k6_needs_bram_9) and (not k4_needs_bram_9)) or ((k1_needs_bram_9) and (not k30_needs_bram_9) and (not k28_needs_bram_9) and (not k26_needs_bram_9) and (not k24_needs_bram_9) and (not k22_needs_bram_9) and (not k20_needs_bram_9) and (not k18_needs_bram_9) and (not k16_needs_bram_9) and (not k14_needs_bram_9) and (not k12_needs_bram_9) and (not k10_needs_bram_9) and (not k8_needs_bram_9) and (not k6_needs_bram_9) and (not k4_needs_bram_9) and (not k2_needs_bram_9));
	bram_21_input_sel(0) <= (k31_needs_bram_10) or ((k29_needs_bram_10) and (not k30_needs_bram_10)) or ((k27_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10)) or ((k25_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10)) or ((k23_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10)) or ((k21_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10)) or ((k19_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10)) or ((k17_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10)) or ((k15_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10)) or ((k13_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10)) or ((k11_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10) and (not k12_needs_bram_10)) or ((k9_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10) and (not k12_needs_bram_10) and (not k10_needs_bram_10)) or ((k7_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10) and (not k12_needs_bram_10) and (not k10_needs_bram_10) and (not k8_needs_bram_10)) or ((k5_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10) and (not k12_needs_bram_10) and (not k10_needs_bram_10) and (not k8_needs_bram_10) and (not k6_needs_bram_10)) or ((k3_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10) and (not k12_needs_bram_10) and (not k10_needs_bram_10) and (not k8_needs_bram_10) and (not k6_needs_bram_10) and (not k4_needs_bram_10)) or ((k1_needs_bram_10) and (not k30_needs_bram_10) and (not k28_needs_bram_10) and (not k26_needs_bram_10) and (not k24_needs_bram_10) and (not k22_needs_bram_10) and (not k20_needs_bram_10) and (not k18_needs_bram_10) and (not k16_needs_bram_10) and (not k14_needs_bram_10) and (not k12_needs_bram_10) and (not k10_needs_bram_10) and (not k8_needs_bram_10) and (not k6_needs_bram_10) and (not k4_needs_bram_10) and (not k2_needs_bram_10));
	bram_23_input_sel(0) <= (k31_needs_bram_11) or ((k29_needs_bram_11) and (not k30_needs_bram_11)) or ((k27_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11)) or ((k25_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11)) or ((k23_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11)) or ((k21_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11)) or ((k19_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11)) or ((k17_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11)) or ((k15_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11)) or ((k13_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11)) or ((k11_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11) and (not k12_needs_bram_11)) or ((k9_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11) and (not k12_needs_bram_11) and (not k10_needs_bram_11)) or ((k7_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11) and (not k12_needs_bram_11) and (not k10_needs_bram_11) and (not k8_needs_bram_11)) or ((k5_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11) and (not k12_needs_bram_11) and (not k10_needs_bram_11) and (not k8_needs_bram_11) and (not k6_needs_bram_11)) or ((k3_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11) and (not k12_needs_bram_11) and (not k10_needs_bram_11) and (not k8_needs_bram_11) and (not k6_needs_bram_11) and (not k4_needs_bram_11)) or ((k1_needs_bram_11) and (not k30_needs_bram_11) and (not k28_needs_bram_11) and (not k26_needs_bram_11) and (not k24_needs_bram_11) and (not k22_needs_bram_11) and (not k20_needs_bram_11) and (not k18_needs_bram_11) and (not k16_needs_bram_11) and (not k14_needs_bram_11) and (not k12_needs_bram_11) and (not k10_needs_bram_11) and (not k8_needs_bram_11) and (not k6_needs_bram_11) and (not k4_needs_bram_11) and (not k2_needs_bram_11));
	bram_25_input_sel(0) <= (k31_needs_bram_12) or ((k29_needs_bram_12) and (not k30_needs_bram_12)) or ((k27_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12)) or ((k25_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12)) or ((k23_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12)) or ((k21_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12)) or ((k19_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12)) or ((k17_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12)) or ((k15_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12)) or ((k13_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12)) or ((k11_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12) and (not k12_needs_bram_12)) or ((k9_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12) and (not k12_needs_bram_12) and (not k10_needs_bram_12)) or ((k7_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12) and (not k12_needs_bram_12) and (not k10_needs_bram_12) and (not k8_needs_bram_12)) or ((k5_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12) and (not k12_needs_bram_12) and (not k10_needs_bram_12) and (not k8_needs_bram_12) and (not k6_needs_bram_12)) or ((k3_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12) and (not k12_needs_bram_12) and (not k10_needs_bram_12) and (not k8_needs_bram_12) and (not k6_needs_bram_12) and (not k4_needs_bram_12)) or ((k1_needs_bram_12) and (not k30_needs_bram_12) and (not k28_needs_bram_12) and (not k26_needs_bram_12) and (not k24_needs_bram_12) and (not k22_needs_bram_12) and (not k20_needs_bram_12) and (not k18_needs_bram_12) and (not k16_needs_bram_12) and (not k14_needs_bram_12) and (not k12_needs_bram_12) and (not k10_needs_bram_12) and (not k8_needs_bram_12) and (not k6_needs_bram_12) and (not k4_needs_bram_12) and (not k2_needs_bram_12));
	bram_27_input_sel(0) <= (k31_needs_bram_13) or ((k29_needs_bram_13) and (not k30_needs_bram_13)) or ((k27_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13)) or ((k25_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13)) or ((k23_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13)) or ((k21_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13)) or ((k19_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13)) or ((k17_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13)) or ((k15_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13)) or ((k13_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13)) or ((k11_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13) and (not k12_needs_bram_13)) or ((k9_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13) and (not k12_needs_bram_13) and (not k10_needs_bram_13)) or ((k7_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13) and (not k12_needs_bram_13) and (not k10_needs_bram_13) and (not k8_needs_bram_13)) or ((k5_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13) and (not k12_needs_bram_13) and (not k10_needs_bram_13) and (not k8_needs_bram_13) and (not k6_needs_bram_13)) or ((k3_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13) and (not k12_needs_bram_13) and (not k10_needs_bram_13) and (not k8_needs_bram_13) and (not k6_needs_bram_13) and (not k4_needs_bram_13)) or ((k1_needs_bram_13) and (not k30_needs_bram_13) and (not k28_needs_bram_13) and (not k26_needs_bram_13) and (not k24_needs_bram_13) and (not k22_needs_bram_13) and (not k20_needs_bram_13) and (not k18_needs_bram_13) and (not k16_needs_bram_13) and (not k14_needs_bram_13) and (not k12_needs_bram_13) and (not k10_needs_bram_13) and (not k8_needs_bram_13) and (not k6_needs_bram_13) and (not k4_needs_bram_13) and (not k2_needs_bram_13));
	bram_29_input_sel(0) <= (k31_needs_bram_14) or ((k29_needs_bram_14) and (not k30_needs_bram_14)) or ((k27_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14)) or ((k25_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14)) or ((k23_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14)) or ((k21_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14)) or ((k19_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14)) or ((k17_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14)) or ((k15_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14)) or ((k13_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14)) or ((k11_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14) and (not k12_needs_bram_14)) or ((k9_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14) and (not k12_needs_bram_14) and (not k10_needs_bram_14)) or ((k7_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14) and (not k12_needs_bram_14) and (not k10_needs_bram_14) and (not k8_needs_bram_14)) or ((k5_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14) and (not k12_needs_bram_14) and (not k10_needs_bram_14) and (not k8_needs_bram_14) and (not k6_needs_bram_14)) or ((k3_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14) and (not k12_needs_bram_14) and (not k10_needs_bram_14) and (not k8_needs_bram_14) and (not k6_needs_bram_14) and (not k4_needs_bram_14)) or ((k1_needs_bram_14) and (not k30_needs_bram_14) and (not k28_needs_bram_14) and (not k26_needs_bram_14) and (not k24_needs_bram_14) and (not k22_needs_bram_14) and (not k20_needs_bram_14) and (not k18_needs_bram_14) and (not k16_needs_bram_14) and (not k14_needs_bram_14) and (not k12_needs_bram_14) and (not k10_needs_bram_14) and (not k8_needs_bram_14) and (not k6_needs_bram_14) and (not k4_needs_bram_14) and (not k2_needs_bram_14));
	bram_31_input_sel(0) <= (k31_needs_bram_15) or ((k29_needs_bram_15) and (not k30_needs_bram_15)) or ((k27_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15)) or ((k25_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15)) or ((k23_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15)) or ((k21_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15)) or ((k19_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15)) or ((k17_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15)) or ((k15_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15)) or ((k13_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15)) or ((k11_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15) and (not k12_needs_bram_15)) or ((k9_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15) and (not k12_needs_bram_15) and (not k10_needs_bram_15)) or ((k7_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15) and (not k12_needs_bram_15) and (not k10_needs_bram_15) and (not k8_needs_bram_15)) or ((k5_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15) and (not k12_needs_bram_15) and (not k10_needs_bram_15) and (not k8_needs_bram_15) and (not k6_needs_bram_15)) or ((k3_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15) and (not k12_needs_bram_15) and (not k10_needs_bram_15) and (not k8_needs_bram_15) and (not k6_needs_bram_15) and (not k4_needs_bram_15)) or ((k1_needs_bram_15) and (not k30_needs_bram_15) and (not k28_needs_bram_15) and (not k26_needs_bram_15) and (not k24_needs_bram_15) and (not k22_needs_bram_15) and (not k20_needs_bram_15) and (not k18_needs_bram_15) and (not k16_needs_bram_15) and (not k14_needs_bram_15) and (not k12_needs_bram_15) and (not k10_needs_bram_15) and (not k8_needs_bram_15) and (not k6_needs_bram_15) and (not k4_needs_bram_15) and (not k2_needs_bram_15));


	addr_0_eq_addr_1 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_1(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_1(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_1(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_1(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_1(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_1(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_1(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_1(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_1(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_1(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_1(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_1(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_1(0))) );

	addr_0_eq_addr_2 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_2(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_2(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_2(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_2(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_2(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_2(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_2(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_2(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_2(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_2(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_2(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_2(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_2(0))) );

	addr_0_eq_addr_3 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_3(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_3(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_3(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_3(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_3(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_3(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_3(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_3(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_3(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_3(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_3(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_3(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_3(0))) );

	addr_0_eq_addr_4 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_4(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_4(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_4(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_4(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_4(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_4(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_4(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_4(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_4(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_4(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_4(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_4(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_4(0))) );

	addr_0_eq_addr_5 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_5(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_5(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_5(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_5(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_5(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_5(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_5(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_5(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_5(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_5(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_5(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_5(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_5(0))) );

	addr_0_eq_addr_6 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_6(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_6(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_6(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_6(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_6(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_6(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_6(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_6(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_6(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_6(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_6(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_6(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_6(0))) );

	addr_0_eq_addr_7 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_7(0))) );

	addr_0_eq_addr_8 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_8(0))) );

	addr_0_eq_addr_9 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_9(0))) );

	addr_0_eq_addr_10 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_10(0))) );

	addr_0_eq_addr_11 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_11(0))) );

	addr_0_eq_addr_12 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_12(0))) );

	addr_0_eq_addr_13 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_13(0))) );

	addr_0_eq_addr_14 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_14(0))) );

	addr_0_eq_addr_15 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_15(0))) );

	addr_0_eq_addr_16 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_16(0))) );

	addr_0_eq_addr_17 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_17(0))) );

	addr_0_eq_addr_18 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_18(0))) );

	addr_0_eq_addr_19 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_19(0))) );

	addr_0_eq_addr_20 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_20(0))) );

	addr_0_eq_addr_21 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_21(0))) );

	addr_0_eq_addr_22 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_22(0))) );

	addr_0_eq_addr_23 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_23(0))) );

	addr_0_eq_addr_24 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_24(0))) );

	addr_0_eq_addr_25 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_25(0))) );

	addr_0_eq_addr_26 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_26(0))) );

	addr_0_eq_addr_27 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_27(0))) );

	addr_0_eq_addr_28 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_28(0))) );

	addr_0_eq_addr_29 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_29(0))) );

	addr_0_eq_addr_30 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_30(0))) );

	addr_0_eq_addr_31 <= ( (to_bit(ADDR_0(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_0(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_0(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_0(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_0(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_0(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_0(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_0(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_0(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_0(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_0(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_0(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_0(0)) xnor to_bit(ADDR_31(0))) );

	addr_1_eq_addr_2 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_2(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_2(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_2(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_2(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_2(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_2(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_2(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_2(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_2(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_2(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_2(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_2(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_2(0))) );

	addr_1_eq_addr_3 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_3(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_3(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_3(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_3(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_3(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_3(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_3(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_3(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_3(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_3(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_3(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_3(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_3(0))) );

	addr_1_eq_addr_4 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_4(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_4(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_4(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_4(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_4(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_4(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_4(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_4(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_4(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_4(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_4(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_4(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_4(0))) );

	addr_1_eq_addr_5 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_5(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_5(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_5(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_5(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_5(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_5(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_5(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_5(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_5(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_5(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_5(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_5(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_5(0))) );

	addr_1_eq_addr_6 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_6(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_6(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_6(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_6(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_6(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_6(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_6(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_6(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_6(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_6(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_6(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_6(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_6(0))) );

	addr_1_eq_addr_7 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_7(0))) );

	addr_1_eq_addr_8 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_8(0))) );

	addr_1_eq_addr_9 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_9(0))) );

	addr_1_eq_addr_10 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_10(0))) );

	addr_1_eq_addr_11 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_11(0))) );

	addr_1_eq_addr_12 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_12(0))) );

	addr_1_eq_addr_13 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_13(0))) );

	addr_1_eq_addr_14 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_14(0))) );

	addr_1_eq_addr_15 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_15(0))) );

	addr_1_eq_addr_16 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_16(0))) );

	addr_1_eq_addr_17 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_17(0))) );

	addr_1_eq_addr_18 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_18(0))) );

	addr_1_eq_addr_19 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_19(0))) );

	addr_1_eq_addr_20 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_20(0))) );

	addr_1_eq_addr_21 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_21(0))) );

	addr_1_eq_addr_22 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_22(0))) );

	addr_1_eq_addr_23 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_23(0))) );

	addr_1_eq_addr_24 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_24(0))) );

	addr_1_eq_addr_25 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_25(0))) );

	addr_1_eq_addr_26 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_26(0))) );

	addr_1_eq_addr_27 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_27(0))) );

	addr_1_eq_addr_28 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_28(0))) );

	addr_1_eq_addr_29 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_29(0))) );

	addr_1_eq_addr_30 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_30(0))) );

	addr_1_eq_addr_31 <= ( (to_bit(ADDR_1(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_1(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_1(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_1(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_1(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_1(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_1(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_1(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_1(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_1(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_1(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_1(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_1(0)) xnor to_bit(ADDR_31(0))) );

	addr_2_eq_addr_3 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_3(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_3(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_3(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_3(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_3(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_3(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_3(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_3(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_3(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_3(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_3(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_3(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_3(0))) );

	addr_2_eq_addr_4 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_4(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_4(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_4(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_4(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_4(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_4(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_4(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_4(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_4(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_4(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_4(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_4(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_4(0))) );

	addr_2_eq_addr_5 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_5(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_5(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_5(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_5(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_5(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_5(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_5(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_5(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_5(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_5(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_5(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_5(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_5(0))) );

	addr_2_eq_addr_6 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_6(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_6(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_6(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_6(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_6(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_6(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_6(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_6(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_6(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_6(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_6(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_6(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_6(0))) );

	addr_2_eq_addr_7 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_7(0))) );

	addr_2_eq_addr_8 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_8(0))) );

	addr_2_eq_addr_9 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_9(0))) );

	addr_2_eq_addr_10 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_10(0))) );

	addr_2_eq_addr_11 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_11(0))) );

	addr_2_eq_addr_12 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_12(0))) );

	addr_2_eq_addr_13 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_13(0))) );

	addr_2_eq_addr_14 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_14(0))) );

	addr_2_eq_addr_15 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_15(0))) );

	addr_2_eq_addr_16 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_16(0))) );

	addr_2_eq_addr_17 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_17(0))) );

	addr_2_eq_addr_18 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_18(0))) );

	addr_2_eq_addr_19 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_19(0))) );

	addr_2_eq_addr_20 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_20(0))) );

	addr_2_eq_addr_21 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_21(0))) );

	addr_2_eq_addr_22 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_22(0))) );

	addr_2_eq_addr_23 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_23(0))) );

	addr_2_eq_addr_24 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_24(0))) );

	addr_2_eq_addr_25 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_25(0))) );

	addr_2_eq_addr_26 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_26(0))) );

	addr_2_eq_addr_27 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_27(0))) );

	addr_2_eq_addr_28 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_28(0))) );

	addr_2_eq_addr_29 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_29(0))) );

	addr_2_eq_addr_30 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_30(0))) );

	addr_2_eq_addr_31 <= ( (to_bit(ADDR_2(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_2(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_2(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_2(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_2(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_2(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_2(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_2(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_2(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_2(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_2(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_2(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_2(0)) xnor to_bit(ADDR_31(0))) );

	addr_3_eq_addr_4 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_4(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_4(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_4(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_4(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_4(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_4(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_4(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_4(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_4(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_4(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_4(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_4(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_4(0))) );

	addr_3_eq_addr_5 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_5(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_5(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_5(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_5(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_5(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_5(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_5(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_5(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_5(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_5(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_5(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_5(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_5(0))) );

	addr_3_eq_addr_6 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_6(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_6(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_6(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_6(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_6(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_6(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_6(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_6(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_6(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_6(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_6(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_6(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_6(0))) );

	addr_3_eq_addr_7 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_7(0))) );

	addr_3_eq_addr_8 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_8(0))) );

	addr_3_eq_addr_9 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_9(0))) );

	addr_3_eq_addr_10 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_10(0))) );

	addr_3_eq_addr_11 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_11(0))) );

	addr_3_eq_addr_12 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_12(0))) );

	addr_3_eq_addr_13 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_13(0))) );

	addr_3_eq_addr_14 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_14(0))) );

	addr_3_eq_addr_15 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_15(0))) );

	addr_3_eq_addr_16 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_16(0))) );

	addr_3_eq_addr_17 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_17(0))) );

	addr_3_eq_addr_18 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_18(0))) );

	addr_3_eq_addr_19 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_19(0))) );

	addr_3_eq_addr_20 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_20(0))) );

	addr_3_eq_addr_21 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_21(0))) );

	addr_3_eq_addr_22 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_22(0))) );

	addr_3_eq_addr_23 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_23(0))) );

	addr_3_eq_addr_24 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_24(0))) );

	addr_3_eq_addr_25 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_25(0))) );

	addr_3_eq_addr_26 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_26(0))) );

	addr_3_eq_addr_27 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_27(0))) );

	addr_3_eq_addr_28 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_28(0))) );

	addr_3_eq_addr_29 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_29(0))) );

	addr_3_eq_addr_30 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_30(0))) );

	addr_3_eq_addr_31 <= ( (to_bit(ADDR_3(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_3(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_3(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_3(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_3(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_3(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_3(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_3(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_3(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_3(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_3(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_3(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_3(0)) xnor to_bit(ADDR_31(0))) );

	addr_4_eq_addr_5 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_5(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_5(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_5(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_5(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_5(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_5(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_5(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_5(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_5(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_5(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_5(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_5(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_5(0))) );

	addr_4_eq_addr_6 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_6(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_6(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_6(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_6(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_6(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_6(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_6(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_6(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_6(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_6(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_6(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_6(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_6(0))) );

	addr_4_eq_addr_7 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_7(0))) );

	addr_4_eq_addr_8 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_8(0))) );

	addr_4_eq_addr_9 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_9(0))) );

	addr_4_eq_addr_10 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_10(0))) );

	addr_4_eq_addr_11 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_11(0))) );

	addr_4_eq_addr_12 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_12(0))) );

	addr_4_eq_addr_13 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_13(0))) );

	addr_4_eq_addr_14 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_14(0))) );

	addr_4_eq_addr_15 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_15(0))) );

	addr_4_eq_addr_16 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_16(0))) );

	addr_4_eq_addr_17 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_17(0))) );

	addr_4_eq_addr_18 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_18(0))) );

	addr_4_eq_addr_19 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_19(0))) );

	addr_4_eq_addr_20 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_20(0))) );

	addr_4_eq_addr_21 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_21(0))) );

	addr_4_eq_addr_22 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_22(0))) );

	addr_4_eq_addr_23 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_23(0))) );

	addr_4_eq_addr_24 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_24(0))) );

	addr_4_eq_addr_25 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_25(0))) );

	addr_4_eq_addr_26 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_26(0))) );

	addr_4_eq_addr_27 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_27(0))) );

	addr_4_eq_addr_28 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_28(0))) );

	addr_4_eq_addr_29 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_29(0))) );

	addr_4_eq_addr_30 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_30(0))) );

	addr_4_eq_addr_31 <= ( (to_bit(ADDR_4(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_4(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_4(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_4(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_4(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_4(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_4(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_4(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_4(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_4(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_4(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_4(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_4(0)) xnor to_bit(ADDR_31(0))) );

	addr_5_eq_addr_6 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_6(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_6(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_6(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_6(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_6(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_6(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_6(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_6(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_6(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_6(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_6(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_6(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_6(0))) );

	addr_5_eq_addr_7 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_7(0))) );

	addr_5_eq_addr_8 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_8(0))) );

	addr_5_eq_addr_9 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_9(0))) );

	addr_5_eq_addr_10 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_10(0))) );

	addr_5_eq_addr_11 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_11(0))) );

	addr_5_eq_addr_12 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_12(0))) );

	addr_5_eq_addr_13 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_13(0))) );

	addr_5_eq_addr_14 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_14(0))) );

	addr_5_eq_addr_15 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_15(0))) );

	addr_5_eq_addr_16 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_16(0))) );

	addr_5_eq_addr_17 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_17(0))) );

	addr_5_eq_addr_18 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_18(0))) );

	addr_5_eq_addr_19 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_19(0))) );

	addr_5_eq_addr_20 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_20(0))) );

	addr_5_eq_addr_21 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_21(0))) );

	addr_5_eq_addr_22 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_22(0))) );

	addr_5_eq_addr_23 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_23(0))) );

	addr_5_eq_addr_24 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_24(0))) );

	addr_5_eq_addr_25 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_25(0))) );

	addr_5_eq_addr_26 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_26(0))) );

	addr_5_eq_addr_27 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_27(0))) );

	addr_5_eq_addr_28 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_28(0))) );

	addr_5_eq_addr_29 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_29(0))) );

	addr_5_eq_addr_30 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_30(0))) );

	addr_5_eq_addr_31 <= ( (to_bit(ADDR_5(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_5(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_5(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_5(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_5(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_5(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_5(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_5(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_5(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_5(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_5(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_5(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_5(0)) xnor to_bit(ADDR_31(0))) );

	addr_6_eq_addr_7 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_7(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_7(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_7(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_7(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_7(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_7(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_7(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_7(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_7(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_7(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_7(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_7(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_7(0))) );

	addr_6_eq_addr_8 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_8(0))) );

	addr_6_eq_addr_9 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_9(0))) );

	addr_6_eq_addr_10 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_10(0))) );

	addr_6_eq_addr_11 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_11(0))) );

	addr_6_eq_addr_12 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_12(0))) );

	addr_6_eq_addr_13 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_13(0))) );

	addr_6_eq_addr_14 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_14(0))) );

	addr_6_eq_addr_15 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_15(0))) );

	addr_6_eq_addr_16 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_16(0))) );

	addr_6_eq_addr_17 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_17(0))) );

	addr_6_eq_addr_18 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_18(0))) );

	addr_6_eq_addr_19 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_19(0))) );

	addr_6_eq_addr_20 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_20(0))) );

	addr_6_eq_addr_21 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_21(0))) );

	addr_6_eq_addr_22 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_22(0))) );

	addr_6_eq_addr_23 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_23(0))) );

	addr_6_eq_addr_24 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_24(0))) );

	addr_6_eq_addr_25 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_25(0))) );

	addr_6_eq_addr_26 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_26(0))) );

	addr_6_eq_addr_27 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_27(0))) );

	addr_6_eq_addr_28 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_28(0))) );

	addr_6_eq_addr_29 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_29(0))) );

	addr_6_eq_addr_30 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_30(0))) );

	addr_6_eq_addr_31 <= ( (to_bit(ADDR_6(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_6(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_6(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_6(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_6(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_6(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_6(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_6(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_6(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_6(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_6(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_6(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_6(0)) xnor to_bit(ADDR_31(0))) );

	addr_7_eq_addr_8 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_8(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_8(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_8(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_8(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_8(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_8(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_8(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_8(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_8(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_8(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_8(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_8(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_8(0))) );

	addr_7_eq_addr_9 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_9(0))) );

	addr_7_eq_addr_10 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_10(0))) );

	addr_7_eq_addr_11 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_11(0))) );

	addr_7_eq_addr_12 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_12(0))) );

	addr_7_eq_addr_13 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_13(0))) );

	addr_7_eq_addr_14 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_14(0))) );

	addr_7_eq_addr_15 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_15(0))) );

	addr_7_eq_addr_16 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_16(0))) );

	addr_7_eq_addr_17 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_17(0))) );

	addr_7_eq_addr_18 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_18(0))) );

	addr_7_eq_addr_19 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_19(0))) );

	addr_7_eq_addr_20 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_20(0))) );

	addr_7_eq_addr_21 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_21(0))) );

	addr_7_eq_addr_22 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_22(0))) );

	addr_7_eq_addr_23 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_23(0))) );

	addr_7_eq_addr_24 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_24(0))) );

	addr_7_eq_addr_25 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_25(0))) );

	addr_7_eq_addr_26 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_26(0))) );

	addr_7_eq_addr_27 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_27(0))) );

	addr_7_eq_addr_28 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_28(0))) );

	addr_7_eq_addr_29 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_29(0))) );

	addr_7_eq_addr_30 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_30(0))) );

	addr_7_eq_addr_31 <= ( (to_bit(ADDR_7(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_7(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_7(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_7(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_7(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_7(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_7(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_7(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_7(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_7(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_7(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_7(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_7(0)) xnor to_bit(ADDR_31(0))) );

	addr_8_eq_addr_9 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_9(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_9(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_9(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_9(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_9(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_9(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_9(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_9(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_9(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_9(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_9(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_9(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_9(0))) );

	addr_8_eq_addr_10 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_10(0))) );

	addr_8_eq_addr_11 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_11(0))) );

	addr_8_eq_addr_12 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_12(0))) );

	addr_8_eq_addr_13 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_13(0))) );

	addr_8_eq_addr_14 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_14(0))) );

	addr_8_eq_addr_15 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_15(0))) );

	addr_8_eq_addr_16 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_16(0))) );

	addr_8_eq_addr_17 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_17(0))) );

	addr_8_eq_addr_18 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_18(0))) );

	addr_8_eq_addr_19 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_19(0))) );

	addr_8_eq_addr_20 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_20(0))) );

	addr_8_eq_addr_21 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_21(0))) );

	addr_8_eq_addr_22 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_22(0))) );

	addr_8_eq_addr_23 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_23(0))) );

	addr_8_eq_addr_24 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_24(0))) );

	addr_8_eq_addr_25 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_25(0))) );

	addr_8_eq_addr_26 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_26(0))) );

	addr_8_eq_addr_27 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_27(0))) );

	addr_8_eq_addr_28 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_28(0))) );

	addr_8_eq_addr_29 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_29(0))) );

	addr_8_eq_addr_30 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_30(0))) );

	addr_8_eq_addr_31 <= ( (to_bit(ADDR_8(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_8(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_8(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_8(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_8(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_8(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_8(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_8(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_8(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_8(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_8(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_8(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_8(0)) xnor to_bit(ADDR_31(0))) );

	addr_9_eq_addr_10 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_10(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_10(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_10(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_10(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_10(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_10(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_10(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_10(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_10(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_10(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_10(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_10(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_10(0))) );

	addr_9_eq_addr_11 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_11(0))) );

	addr_9_eq_addr_12 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_12(0))) );

	addr_9_eq_addr_13 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_13(0))) );

	addr_9_eq_addr_14 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_14(0))) );

	addr_9_eq_addr_15 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_15(0))) );

	addr_9_eq_addr_16 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_16(0))) );

	addr_9_eq_addr_17 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_17(0))) );

	addr_9_eq_addr_18 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_18(0))) );

	addr_9_eq_addr_19 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_19(0))) );

	addr_9_eq_addr_20 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_20(0))) );

	addr_9_eq_addr_21 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_21(0))) );

	addr_9_eq_addr_22 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_22(0))) );

	addr_9_eq_addr_23 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_23(0))) );

	addr_9_eq_addr_24 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_24(0))) );

	addr_9_eq_addr_25 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_25(0))) );

	addr_9_eq_addr_26 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_26(0))) );

	addr_9_eq_addr_27 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_27(0))) );

	addr_9_eq_addr_28 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_28(0))) );

	addr_9_eq_addr_29 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_29(0))) );

	addr_9_eq_addr_30 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_30(0))) );

	addr_9_eq_addr_31 <= ( (to_bit(ADDR_9(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_9(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_9(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_9(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_9(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_9(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_9(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_9(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_9(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_9(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_9(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_9(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_9(0)) xnor to_bit(ADDR_31(0))) );

	addr_10_eq_addr_11 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_11(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_11(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_11(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_11(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_11(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_11(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_11(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_11(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_11(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_11(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_11(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_11(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_11(0))) );

	addr_10_eq_addr_12 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_12(0))) );

	addr_10_eq_addr_13 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_13(0))) );

	addr_10_eq_addr_14 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_14(0))) );

	addr_10_eq_addr_15 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_15(0))) );

	addr_10_eq_addr_16 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_16(0))) );

	addr_10_eq_addr_17 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_17(0))) );

	addr_10_eq_addr_18 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_18(0))) );

	addr_10_eq_addr_19 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_19(0))) );

	addr_10_eq_addr_20 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_20(0))) );

	addr_10_eq_addr_21 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_21(0))) );

	addr_10_eq_addr_22 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_22(0))) );

	addr_10_eq_addr_23 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_23(0))) );

	addr_10_eq_addr_24 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_24(0))) );

	addr_10_eq_addr_25 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_25(0))) );

	addr_10_eq_addr_26 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_26(0))) );

	addr_10_eq_addr_27 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_27(0))) );

	addr_10_eq_addr_28 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_28(0))) );

	addr_10_eq_addr_29 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_29(0))) );

	addr_10_eq_addr_30 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_30(0))) );

	addr_10_eq_addr_31 <= ( (to_bit(ADDR_10(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_10(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_10(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_10(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_10(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_10(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_10(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_10(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_10(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_10(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_10(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_10(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_10(0)) xnor to_bit(ADDR_31(0))) );

	addr_11_eq_addr_12 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_12(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_12(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_12(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_12(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_12(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_12(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_12(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_12(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_12(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_12(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_12(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_12(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_12(0))) );

	addr_11_eq_addr_13 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_13(0))) );

	addr_11_eq_addr_14 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_14(0))) );

	addr_11_eq_addr_15 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_15(0))) );

	addr_11_eq_addr_16 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_16(0))) );

	addr_11_eq_addr_17 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_17(0))) );

	addr_11_eq_addr_18 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_18(0))) );

	addr_11_eq_addr_19 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_19(0))) );

	addr_11_eq_addr_20 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_20(0))) );

	addr_11_eq_addr_21 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_21(0))) );

	addr_11_eq_addr_22 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_22(0))) );

	addr_11_eq_addr_23 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_23(0))) );

	addr_11_eq_addr_24 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_24(0))) );

	addr_11_eq_addr_25 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_25(0))) );

	addr_11_eq_addr_26 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_26(0))) );

	addr_11_eq_addr_27 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_27(0))) );

	addr_11_eq_addr_28 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_28(0))) );

	addr_11_eq_addr_29 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_29(0))) );

	addr_11_eq_addr_30 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_30(0))) );

	addr_11_eq_addr_31 <= ( (to_bit(ADDR_11(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_11(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_11(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_11(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_11(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_11(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_11(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_11(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_11(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_11(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_11(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_11(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_11(0)) xnor to_bit(ADDR_31(0))) );

	addr_12_eq_addr_13 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_13(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_13(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_13(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_13(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_13(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_13(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_13(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_13(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_13(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_13(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_13(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_13(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_13(0))) );

	addr_12_eq_addr_14 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_14(0))) );

	addr_12_eq_addr_15 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_15(0))) );

	addr_12_eq_addr_16 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_16(0))) );

	addr_12_eq_addr_17 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_17(0))) );

	addr_12_eq_addr_18 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_18(0))) );

	addr_12_eq_addr_19 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_19(0))) );

	addr_12_eq_addr_20 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_20(0))) );

	addr_12_eq_addr_21 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_21(0))) );

	addr_12_eq_addr_22 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_22(0))) );

	addr_12_eq_addr_23 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_23(0))) );

	addr_12_eq_addr_24 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_24(0))) );

	addr_12_eq_addr_25 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_25(0))) );

	addr_12_eq_addr_26 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_26(0))) );

	addr_12_eq_addr_27 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_27(0))) );

	addr_12_eq_addr_28 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_28(0))) );

	addr_12_eq_addr_29 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_29(0))) );

	addr_12_eq_addr_30 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_30(0))) );

	addr_12_eq_addr_31 <= ( (to_bit(ADDR_12(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_12(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_12(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_12(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_12(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_12(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_12(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_12(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_12(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_12(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_12(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_12(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_12(0)) xnor to_bit(ADDR_31(0))) );

	addr_13_eq_addr_14 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_14(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_14(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_14(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_14(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_14(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_14(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_14(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_14(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_14(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_14(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_14(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_14(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_14(0))) );

	addr_13_eq_addr_15 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_15(0))) );

	addr_13_eq_addr_16 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_16(0))) );

	addr_13_eq_addr_17 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_17(0))) );

	addr_13_eq_addr_18 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_18(0))) );

	addr_13_eq_addr_19 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_19(0))) );

	addr_13_eq_addr_20 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_20(0))) );

	addr_13_eq_addr_21 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_21(0))) );

	addr_13_eq_addr_22 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_22(0))) );

	addr_13_eq_addr_23 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_23(0))) );

	addr_13_eq_addr_24 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_24(0))) );

	addr_13_eq_addr_25 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_25(0))) );

	addr_13_eq_addr_26 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_26(0))) );

	addr_13_eq_addr_27 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_27(0))) );

	addr_13_eq_addr_28 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_28(0))) );

	addr_13_eq_addr_29 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_29(0))) );

	addr_13_eq_addr_30 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_30(0))) );

	addr_13_eq_addr_31 <= ( (to_bit(ADDR_13(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_13(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_13(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_13(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_13(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_13(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_13(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_13(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_13(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_13(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_13(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_13(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_13(0)) xnor to_bit(ADDR_31(0))) );

	addr_14_eq_addr_15 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_15(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_15(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_15(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_15(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_15(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_15(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_15(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_15(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_15(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_15(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_15(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_15(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_15(0))) );

	addr_14_eq_addr_16 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_16(0))) );

	addr_14_eq_addr_17 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_17(0))) );

	addr_14_eq_addr_18 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_18(0))) );

	addr_14_eq_addr_19 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_19(0))) );

	addr_14_eq_addr_20 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_20(0))) );

	addr_14_eq_addr_21 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_21(0))) );

	addr_14_eq_addr_22 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_22(0))) );

	addr_14_eq_addr_23 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_23(0))) );

	addr_14_eq_addr_24 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_24(0))) );

	addr_14_eq_addr_25 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_25(0))) );

	addr_14_eq_addr_26 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_26(0))) );

	addr_14_eq_addr_27 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_27(0))) );

	addr_14_eq_addr_28 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_28(0))) );

	addr_14_eq_addr_29 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_29(0))) );

	addr_14_eq_addr_30 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_30(0))) );

	addr_14_eq_addr_31 <= ( (to_bit(ADDR_14(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_14(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_14(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_14(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_14(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_14(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_14(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_14(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_14(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_14(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_14(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_14(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_14(0)) xnor to_bit(ADDR_31(0))) );

	addr_15_eq_addr_16 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_16(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_16(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_16(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_16(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_16(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_16(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_16(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_16(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_16(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_16(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_16(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_16(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_16(0))) );

	addr_15_eq_addr_17 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_17(0))) );

	addr_15_eq_addr_18 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_18(0))) );

	addr_15_eq_addr_19 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_19(0))) );

	addr_15_eq_addr_20 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_20(0))) );

	addr_15_eq_addr_21 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_21(0))) );

	addr_15_eq_addr_22 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_22(0))) );

	addr_15_eq_addr_23 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_23(0))) );

	addr_15_eq_addr_24 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_24(0))) );

	addr_15_eq_addr_25 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_25(0))) );

	addr_15_eq_addr_26 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_26(0))) );

	addr_15_eq_addr_27 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_27(0))) );

	addr_15_eq_addr_28 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_28(0))) );

	addr_15_eq_addr_29 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_29(0))) );

	addr_15_eq_addr_30 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_30(0))) );

	addr_15_eq_addr_31 <= ( (to_bit(ADDR_15(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_15(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_15(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_15(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_15(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_15(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_15(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_15(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_15(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_15(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_15(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_15(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_15(0)) xnor to_bit(ADDR_31(0))) );

	addr_16_eq_addr_17 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_17(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_17(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_17(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_17(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_17(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_17(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_17(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_17(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_17(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_17(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_17(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_17(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_17(0))) );

	addr_16_eq_addr_18 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_18(0))) );

	addr_16_eq_addr_19 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_19(0))) );

	addr_16_eq_addr_20 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_20(0))) );

	addr_16_eq_addr_21 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_21(0))) );

	addr_16_eq_addr_22 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_22(0))) );

	addr_16_eq_addr_23 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_23(0))) );

	addr_16_eq_addr_24 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_24(0))) );

	addr_16_eq_addr_25 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_25(0))) );

	addr_16_eq_addr_26 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_26(0))) );

	addr_16_eq_addr_27 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_27(0))) );

	addr_16_eq_addr_28 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_28(0))) );

	addr_16_eq_addr_29 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_29(0))) );

	addr_16_eq_addr_30 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_30(0))) );

	addr_16_eq_addr_31 <= ( (to_bit(ADDR_16(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_16(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_16(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_16(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_16(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_16(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_16(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_16(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_16(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_16(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_16(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_16(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_16(0)) xnor to_bit(ADDR_31(0))) );

	addr_17_eq_addr_18 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_18(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_18(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_18(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_18(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_18(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_18(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_18(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_18(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_18(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_18(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_18(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_18(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_18(0))) );

	addr_17_eq_addr_19 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_19(0))) );

	addr_17_eq_addr_20 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_20(0))) );

	addr_17_eq_addr_21 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_21(0))) );

	addr_17_eq_addr_22 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_22(0))) );

	addr_17_eq_addr_23 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_23(0))) );

	addr_17_eq_addr_24 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_24(0))) );

	addr_17_eq_addr_25 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_25(0))) );

	addr_17_eq_addr_26 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_26(0))) );

	addr_17_eq_addr_27 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_27(0))) );

	addr_17_eq_addr_28 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_28(0))) );

	addr_17_eq_addr_29 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_29(0))) );

	addr_17_eq_addr_30 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_30(0))) );

	addr_17_eq_addr_31 <= ( (to_bit(ADDR_17(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_17(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_17(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_17(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_17(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_17(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_17(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_17(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_17(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_17(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_17(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_17(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_17(0)) xnor to_bit(ADDR_31(0))) );

	addr_18_eq_addr_19 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_19(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_19(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_19(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_19(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_19(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_19(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_19(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_19(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_19(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_19(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_19(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_19(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_19(0))) );

	addr_18_eq_addr_20 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_20(0))) );

	addr_18_eq_addr_21 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_21(0))) );

	addr_18_eq_addr_22 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_22(0))) );

	addr_18_eq_addr_23 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_23(0))) );

	addr_18_eq_addr_24 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_24(0))) );

	addr_18_eq_addr_25 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_25(0))) );

	addr_18_eq_addr_26 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_26(0))) );

	addr_18_eq_addr_27 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_27(0))) );

	addr_18_eq_addr_28 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_28(0))) );

	addr_18_eq_addr_29 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_29(0))) );

	addr_18_eq_addr_30 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_30(0))) );

	addr_18_eq_addr_31 <= ( (to_bit(ADDR_18(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_18(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_18(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_18(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_18(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_18(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_18(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_18(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_18(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_18(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_18(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_18(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_18(0)) xnor to_bit(ADDR_31(0))) );

	addr_19_eq_addr_20 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_20(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_20(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_20(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_20(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_20(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_20(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_20(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_20(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_20(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_20(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_20(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_20(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_20(0))) );

	addr_19_eq_addr_21 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_21(0))) );

	addr_19_eq_addr_22 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_22(0))) );

	addr_19_eq_addr_23 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_23(0))) );

	addr_19_eq_addr_24 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_24(0))) );

	addr_19_eq_addr_25 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_25(0))) );

	addr_19_eq_addr_26 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_26(0))) );

	addr_19_eq_addr_27 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_27(0))) );

	addr_19_eq_addr_28 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_28(0))) );

	addr_19_eq_addr_29 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_29(0))) );

	addr_19_eq_addr_30 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_30(0))) );

	addr_19_eq_addr_31 <= ( (to_bit(ADDR_19(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_19(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_19(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_19(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_19(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_19(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_19(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_19(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_19(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_19(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_19(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_19(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_19(0)) xnor to_bit(ADDR_31(0))) );

	addr_20_eq_addr_21 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_21(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_21(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_21(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_21(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_21(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_21(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_21(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_21(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_21(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_21(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_21(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_21(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_21(0))) );

	addr_20_eq_addr_22 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_22(0))) );

	addr_20_eq_addr_23 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_23(0))) );

	addr_20_eq_addr_24 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_24(0))) );

	addr_20_eq_addr_25 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_25(0))) );

	addr_20_eq_addr_26 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_26(0))) );

	addr_20_eq_addr_27 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_27(0))) );

	addr_20_eq_addr_28 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_28(0))) );

	addr_20_eq_addr_29 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_29(0))) );

	addr_20_eq_addr_30 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_30(0))) );

	addr_20_eq_addr_31 <= ( (to_bit(ADDR_20(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_20(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_20(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_20(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_20(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_20(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_20(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_20(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_20(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_20(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_20(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_20(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_20(0)) xnor to_bit(ADDR_31(0))) );

	addr_21_eq_addr_22 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_22(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_22(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_22(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_22(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_22(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_22(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_22(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_22(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_22(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_22(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_22(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_22(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_22(0))) );

	addr_21_eq_addr_23 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_23(0))) );

	addr_21_eq_addr_24 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_24(0))) );

	addr_21_eq_addr_25 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_25(0))) );

	addr_21_eq_addr_26 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_26(0))) );

	addr_21_eq_addr_27 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_27(0))) );

	addr_21_eq_addr_28 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_28(0))) );

	addr_21_eq_addr_29 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_29(0))) );

	addr_21_eq_addr_30 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_30(0))) );

	addr_21_eq_addr_31 <= ( (to_bit(ADDR_21(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_21(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_21(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_21(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_21(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_21(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_21(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_21(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_21(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_21(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_21(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_21(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_21(0)) xnor to_bit(ADDR_31(0))) );

	addr_22_eq_addr_23 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_23(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_23(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_23(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_23(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_23(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_23(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_23(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_23(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_23(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_23(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_23(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_23(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_23(0))) );

	addr_22_eq_addr_24 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_24(0))) );

	addr_22_eq_addr_25 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_25(0))) );

	addr_22_eq_addr_26 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_26(0))) );

	addr_22_eq_addr_27 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_27(0))) );

	addr_22_eq_addr_28 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_28(0))) );

	addr_22_eq_addr_29 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_29(0))) );

	addr_22_eq_addr_30 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_30(0))) );

	addr_22_eq_addr_31 <= ( (to_bit(ADDR_22(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_22(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_22(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_22(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_22(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_22(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_22(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_22(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_22(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_22(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_22(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_22(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_22(0)) xnor to_bit(ADDR_31(0))) );

	addr_23_eq_addr_24 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_24(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_24(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_24(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_24(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_24(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_24(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_24(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_24(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_24(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_24(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_24(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_24(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_24(0))) );

	addr_23_eq_addr_25 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_25(0))) );

	addr_23_eq_addr_26 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_26(0))) );

	addr_23_eq_addr_27 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_27(0))) );

	addr_23_eq_addr_28 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_28(0))) );

	addr_23_eq_addr_29 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_29(0))) );

	addr_23_eq_addr_30 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_30(0))) );

	addr_23_eq_addr_31 <= ( (to_bit(ADDR_23(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_23(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_23(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_23(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_23(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_23(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_23(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_23(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_23(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_23(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_23(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_23(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_23(0)) xnor to_bit(ADDR_31(0))) );

	addr_24_eq_addr_25 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_25(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_25(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_25(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_25(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_25(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_25(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_25(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_25(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_25(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_25(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_25(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_25(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_25(0))) );

	addr_24_eq_addr_26 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_26(0))) );

	addr_24_eq_addr_27 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_27(0))) );

	addr_24_eq_addr_28 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_28(0))) );

	addr_24_eq_addr_29 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_29(0))) );

	addr_24_eq_addr_30 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_30(0))) );

	addr_24_eq_addr_31 <= ( (to_bit(ADDR_24(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_24(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_24(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_24(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_24(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_24(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_24(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_24(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_24(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_24(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_24(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_24(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_24(0)) xnor to_bit(ADDR_31(0))) );

	addr_25_eq_addr_26 <= ( (to_bit(ADDR_25(12)) xnor to_bit(ADDR_26(12))) and
	                      (to_bit(ADDR_25(11)) xnor to_bit(ADDR_26(11))) and
	                      (to_bit(ADDR_25(10)) xnor to_bit(ADDR_26(10))) and
	                      (to_bit(ADDR_25(9)) xnor to_bit(ADDR_26(9))) and
	                      (to_bit(ADDR_25(8)) xnor to_bit(ADDR_26(8))) and
	                      (to_bit(ADDR_25(7)) xnor to_bit(ADDR_26(7))) and
	                      (to_bit(ADDR_25(6)) xnor to_bit(ADDR_26(6))) and
	                      (to_bit(ADDR_25(5)) xnor to_bit(ADDR_26(5))) and
	                      (to_bit(ADDR_25(4)) xnor to_bit(ADDR_26(4))) and
	                      (to_bit(ADDR_25(3)) xnor to_bit(ADDR_26(3))) and
	                      (to_bit(ADDR_25(2)) xnor to_bit(ADDR_26(2))) and
	                      (to_bit(ADDR_25(1)) xnor to_bit(ADDR_26(1))) and
	                      (to_bit(ADDR_25(0)) xnor to_bit(ADDR_26(0))) );

	addr_25_eq_addr_27 <= ( (to_bit(ADDR_25(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_25(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_25(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_25(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_25(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_25(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_25(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_25(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_25(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_25(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_25(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_25(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_25(0)) xnor to_bit(ADDR_27(0))) );

	addr_25_eq_addr_28 <= ( (to_bit(ADDR_25(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_25(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_25(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_25(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_25(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_25(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_25(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_25(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_25(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_25(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_25(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_25(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_25(0)) xnor to_bit(ADDR_28(0))) );

	addr_25_eq_addr_29 <= ( (to_bit(ADDR_25(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_25(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_25(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_25(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_25(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_25(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_25(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_25(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_25(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_25(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_25(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_25(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_25(0)) xnor to_bit(ADDR_29(0))) );

	addr_25_eq_addr_30 <= ( (to_bit(ADDR_25(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_25(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_25(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_25(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_25(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_25(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_25(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_25(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_25(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_25(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_25(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_25(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_25(0)) xnor to_bit(ADDR_30(0))) );

	addr_25_eq_addr_31 <= ( (to_bit(ADDR_25(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_25(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_25(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_25(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_25(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_25(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_25(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_25(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_25(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_25(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_25(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_25(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_25(0)) xnor to_bit(ADDR_31(0))) );

	addr_26_eq_addr_27 <= ( (to_bit(ADDR_26(12)) xnor to_bit(ADDR_27(12))) and
	                      (to_bit(ADDR_26(11)) xnor to_bit(ADDR_27(11))) and
	                      (to_bit(ADDR_26(10)) xnor to_bit(ADDR_27(10))) and
	                      (to_bit(ADDR_26(9)) xnor to_bit(ADDR_27(9))) and
	                      (to_bit(ADDR_26(8)) xnor to_bit(ADDR_27(8))) and
	                      (to_bit(ADDR_26(7)) xnor to_bit(ADDR_27(7))) and
	                      (to_bit(ADDR_26(6)) xnor to_bit(ADDR_27(6))) and
	                      (to_bit(ADDR_26(5)) xnor to_bit(ADDR_27(5))) and
	                      (to_bit(ADDR_26(4)) xnor to_bit(ADDR_27(4))) and
	                      (to_bit(ADDR_26(3)) xnor to_bit(ADDR_27(3))) and
	                      (to_bit(ADDR_26(2)) xnor to_bit(ADDR_27(2))) and
	                      (to_bit(ADDR_26(1)) xnor to_bit(ADDR_27(1))) and
	                      (to_bit(ADDR_26(0)) xnor to_bit(ADDR_27(0))) );

	addr_26_eq_addr_28 <= ( (to_bit(ADDR_26(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_26(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_26(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_26(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_26(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_26(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_26(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_26(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_26(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_26(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_26(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_26(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_26(0)) xnor to_bit(ADDR_28(0))) );

	addr_26_eq_addr_29 <= ( (to_bit(ADDR_26(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_26(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_26(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_26(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_26(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_26(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_26(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_26(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_26(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_26(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_26(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_26(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_26(0)) xnor to_bit(ADDR_29(0))) );

	addr_26_eq_addr_30 <= ( (to_bit(ADDR_26(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_26(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_26(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_26(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_26(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_26(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_26(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_26(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_26(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_26(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_26(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_26(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_26(0)) xnor to_bit(ADDR_30(0))) );

	addr_26_eq_addr_31 <= ( (to_bit(ADDR_26(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_26(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_26(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_26(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_26(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_26(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_26(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_26(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_26(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_26(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_26(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_26(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_26(0)) xnor to_bit(ADDR_31(0))) );

	addr_27_eq_addr_28 <= ( (to_bit(ADDR_27(12)) xnor to_bit(ADDR_28(12))) and
	                      (to_bit(ADDR_27(11)) xnor to_bit(ADDR_28(11))) and
	                      (to_bit(ADDR_27(10)) xnor to_bit(ADDR_28(10))) and
	                      (to_bit(ADDR_27(9)) xnor to_bit(ADDR_28(9))) and
	                      (to_bit(ADDR_27(8)) xnor to_bit(ADDR_28(8))) and
	                      (to_bit(ADDR_27(7)) xnor to_bit(ADDR_28(7))) and
	                      (to_bit(ADDR_27(6)) xnor to_bit(ADDR_28(6))) and
	                      (to_bit(ADDR_27(5)) xnor to_bit(ADDR_28(5))) and
	                      (to_bit(ADDR_27(4)) xnor to_bit(ADDR_28(4))) and
	                      (to_bit(ADDR_27(3)) xnor to_bit(ADDR_28(3))) and
	                      (to_bit(ADDR_27(2)) xnor to_bit(ADDR_28(2))) and
	                      (to_bit(ADDR_27(1)) xnor to_bit(ADDR_28(1))) and
	                      (to_bit(ADDR_27(0)) xnor to_bit(ADDR_28(0))) );

	addr_27_eq_addr_29 <= ( (to_bit(ADDR_27(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_27(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_27(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_27(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_27(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_27(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_27(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_27(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_27(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_27(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_27(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_27(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_27(0)) xnor to_bit(ADDR_29(0))) );

	addr_27_eq_addr_30 <= ( (to_bit(ADDR_27(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_27(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_27(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_27(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_27(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_27(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_27(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_27(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_27(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_27(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_27(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_27(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_27(0)) xnor to_bit(ADDR_30(0))) );

	addr_27_eq_addr_31 <= ( (to_bit(ADDR_27(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_27(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_27(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_27(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_27(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_27(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_27(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_27(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_27(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_27(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_27(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_27(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_27(0)) xnor to_bit(ADDR_31(0))) );

	addr_28_eq_addr_29 <= ( (to_bit(ADDR_28(12)) xnor to_bit(ADDR_29(12))) and
	                      (to_bit(ADDR_28(11)) xnor to_bit(ADDR_29(11))) and
	                      (to_bit(ADDR_28(10)) xnor to_bit(ADDR_29(10))) and
	                      (to_bit(ADDR_28(9)) xnor to_bit(ADDR_29(9))) and
	                      (to_bit(ADDR_28(8)) xnor to_bit(ADDR_29(8))) and
	                      (to_bit(ADDR_28(7)) xnor to_bit(ADDR_29(7))) and
	                      (to_bit(ADDR_28(6)) xnor to_bit(ADDR_29(6))) and
	                      (to_bit(ADDR_28(5)) xnor to_bit(ADDR_29(5))) and
	                      (to_bit(ADDR_28(4)) xnor to_bit(ADDR_29(4))) and
	                      (to_bit(ADDR_28(3)) xnor to_bit(ADDR_29(3))) and
	                      (to_bit(ADDR_28(2)) xnor to_bit(ADDR_29(2))) and
	                      (to_bit(ADDR_28(1)) xnor to_bit(ADDR_29(1))) and
	                      (to_bit(ADDR_28(0)) xnor to_bit(ADDR_29(0))) );

	addr_28_eq_addr_30 <= ( (to_bit(ADDR_28(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_28(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_28(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_28(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_28(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_28(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_28(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_28(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_28(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_28(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_28(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_28(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_28(0)) xnor to_bit(ADDR_30(0))) );

	addr_28_eq_addr_31 <= ( (to_bit(ADDR_28(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_28(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_28(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_28(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_28(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_28(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_28(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_28(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_28(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_28(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_28(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_28(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_28(0)) xnor to_bit(ADDR_31(0))) );

	addr_29_eq_addr_30 <= ( (to_bit(ADDR_29(12)) xnor to_bit(ADDR_30(12))) and
	                      (to_bit(ADDR_29(11)) xnor to_bit(ADDR_30(11))) and
	                      (to_bit(ADDR_29(10)) xnor to_bit(ADDR_30(10))) and
	                      (to_bit(ADDR_29(9)) xnor to_bit(ADDR_30(9))) and
	                      (to_bit(ADDR_29(8)) xnor to_bit(ADDR_30(8))) and
	                      (to_bit(ADDR_29(7)) xnor to_bit(ADDR_30(7))) and
	                      (to_bit(ADDR_29(6)) xnor to_bit(ADDR_30(6))) and
	                      (to_bit(ADDR_29(5)) xnor to_bit(ADDR_30(5))) and
	                      (to_bit(ADDR_29(4)) xnor to_bit(ADDR_30(4))) and
	                      (to_bit(ADDR_29(3)) xnor to_bit(ADDR_30(3))) and
	                      (to_bit(ADDR_29(2)) xnor to_bit(ADDR_30(2))) and
	                      (to_bit(ADDR_29(1)) xnor to_bit(ADDR_30(1))) and
	                      (to_bit(ADDR_29(0)) xnor to_bit(ADDR_30(0))) );

	addr_29_eq_addr_31 <= ( (to_bit(ADDR_29(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_29(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_29(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_29(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_29(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_29(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_29(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_29(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_29(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_29(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_29(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_29(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_29(0)) xnor to_bit(ADDR_31(0))) );

	addr_30_eq_addr_31 <= ( (to_bit(ADDR_30(12)) xnor to_bit(ADDR_31(12))) and
	                      (to_bit(ADDR_30(11)) xnor to_bit(ADDR_31(11))) and
	                      (to_bit(ADDR_30(10)) xnor to_bit(ADDR_31(10))) and
	                      (to_bit(ADDR_30(9)) xnor to_bit(ADDR_31(9))) and
	                      (to_bit(ADDR_30(8)) xnor to_bit(ADDR_31(8))) and
	                      (to_bit(ADDR_30(7)) xnor to_bit(ADDR_31(7))) and
	                      (to_bit(ADDR_30(6)) xnor to_bit(ADDR_31(6))) and
	                      (to_bit(ADDR_30(5)) xnor to_bit(ADDR_31(5))) and
	                      (to_bit(ADDR_30(4)) xnor to_bit(ADDR_31(4))) and
	                      (to_bit(ADDR_30(3)) xnor to_bit(ADDR_31(3))) and
	                      (to_bit(ADDR_30(2)) xnor to_bit(ADDR_31(2))) and
	                      (to_bit(ADDR_30(1)) xnor to_bit(ADDR_31(1))) and
	                      (to_bit(ADDR_30(0)) xnor to_bit(ADDR_31(0))) );


	k0_being_served <= to_bit(REQ_0);

	k1_being_served <= to_bit(REQ_1) and (
	                       ( not k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and not k1_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and     k1_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k1_needs_attention) );

	k2_being_served <= to_bit(REQ_2) and (
	                       ( not k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and not k2_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and     k2_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k2_needs_attention) );

	k3_being_served <= to_bit(REQ_3) and (
	                       ( not k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and not k3_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and     k3_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k3_needs_attention) );

	k4_being_served <= to_bit(REQ_4) and (
	                       ( not k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and not k4_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and     k4_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k4_needs_attention) );

	k5_being_served <= to_bit(REQ_5) and (
	                       ( not k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and not k5_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and     k5_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k5_needs_attention) );

	k6_being_served <= to_bit(REQ_6) and (
	                       ( not k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and not k6_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and     k6_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k6_needs_attention) );

	k7_being_served <= to_bit(REQ_7) and (
	                       ( not k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and not k7_output_sel(0) and ( ( not bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and     k7_output_sel(0) and ( ( not bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k7_needs_attention) );

	k8_being_served <= to_bit(REQ_8) and (
	                       ( not k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and not k8_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and     k8_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k8_needs_attention) );

	k9_being_served <= to_bit(REQ_9) and (
	                       ( not k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and not k9_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and     k9_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k9_needs_attention) );

	k10_being_served <= to_bit(REQ_10) and (
	                       ( not k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and not k10_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and     k10_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k10_needs_attention) );

	k11_being_served <= to_bit(REQ_11) and (
	                       ( not k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and not k11_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and     k11_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k11_needs_attention) );

	k12_being_served <= to_bit(REQ_12) and (
	                       ( not k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and not k12_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and     k12_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k12_needs_attention) );

	k13_being_served <= to_bit(REQ_13) and (
	                       ( not k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and not k13_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and     k13_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k13_needs_attention) );

	k14_being_served <= to_bit(REQ_14) and (
	                       ( not k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and not k14_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and     k14_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k14_needs_attention) );

	k15_being_served <= to_bit(REQ_15) and (
	                       ( not k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             ( not bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             ( not bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             ( not bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             ( not bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             ( not bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             ( not bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             ( not bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             ( not bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             ( not bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             ( not bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             ( not bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             ( not bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             ( not bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             ( not bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and not k15_output_sel(0) and ( ( not bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             ( not bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and     k15_output_sel(0) and ( ( not bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             ( not bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k15_needs_attention) );

	k16_being_served <= to_bit(REQ_16) and (
	                       ( not k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and not k16_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and     k16_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k16_needs_attention) );

	k17_being_served <= to_bit(REQ_17) and (
	                       ( not k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and not k17_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and     k17_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k17_needs_attention) );

	k18_being_served <= to_bit(REQ_18) and (
	                       ( not k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and not k18_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and     k18_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k18_needs_attention) );

	k19_being_served <= to_bit(REQ_19) and (
	                       ( not k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and not k19_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and     k19_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k19_needs_attention) );

	k20_being_served <= to_bit(REQ_20) and (
	                       ( not k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and not k20_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and     k20_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k20_needs_attention) );

	k21_being_served <= to_bit(REQ_21) and (
	                       ( not k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and not k21_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and     k21_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k21_needs_attention) );

	k22_being_served <= to_bit(REQ_22) and (
	                       ( not k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and not k22_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and     k22_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k22_needs_attention) );

	k23_being_served <= to_bit(REQ_23) and (
	                       ( not k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_0_input_sel(4) and not bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and not bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_2_input_sel(4) and not bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and not bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_4_input_sel(4) and not bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and not bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_6_input_sel(4) and not bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and not bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_8_input_sel(4) and not bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and not bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_10_input_sel(4) and not bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and not bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_12_input_sel(4) and not bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and not bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_14_input_sel(4) and not bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and not bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_16_input_sel(4) and not bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and not bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_18_input_sel(4) and not bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and not bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_20_input_sel(4) and not bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and not bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_22_input_sel(4) and not bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and not bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_24_input_sel(4) and not bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and not bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_26_input_sel(4) and not bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and not bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and not k23_output_sel(0) and ( (     bram_28_input_sel(4) and not bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and not bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and     k23_output_sel(0) and ( (     bram_30_input_sel(4) and not bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and not bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k23_needs_attention) );

	k24_being_served <= to_bit(REQ_24) and (
	                       ( not k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and not k24_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and     k24_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k24_needs_attention) );

	k25_being_served <= to_bit(REQ_25) and (
	                       ( not k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and not k25_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and     k25_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k25_needs_attention) );

	k26_being_served <= to_bit(REQ_26) and (
	                       ( not k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and not k26_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and     k26_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k26_needs_attention) );

	k27_being_served <= to_bit(REQ_27) and (
	                       ( not k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and not bram_0_input_sel(2) and     bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and not bram_1_input_sel(2) and     bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and not bram_2_input_sel(2) and     bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and not bram_3_input_sel(2) and     bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and not bram_4_input_sel(2) and     bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and not bram_5_input_sel(2) and     bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and not bram_6_input_sel(2) and     bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and not bram_7_input_sel(2) and     bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and not bram_8_input_sel(2) and     bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and not bram_9_input_sel(2) and     bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and not bram_10_input_sel(2) and     bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and not bram_11_input_sel(2) and     bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and not bram_12_input_sel(2) and     bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and not bram_13_input_sel(2) and     bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and not bram_14_input_sel(2) and     bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and not bram_15_input_sel(2) and     bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and not bram_16_input_sel(2) and     bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and not bram_17_input_sel(2) and     bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and not bram_18_input_sel(2) and     bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and not bram_19_input_sel(2) and     bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and not bram_20_input_sel(2) and     bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and not bram_21_input_sel(2) and     bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and not bram_22_input_sel(2) and     bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and not bram_23_input_sel(2) and     bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and not bram_24_input_sel(2) and     bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and not bram_25_input_sel(2) and     bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and not bram_26_input_sel(2) and     bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and not bram_27_input_sel(2) and     bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and not k27_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and not bram_28_input_sel(2) and     bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and not bram_29_input_sel(2) and     bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and     k27_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and not bram_30_input_sel(2) and     bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and not bram_31_input_sel(2) and     bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k27_needs_attention) );

	k28_being_served <= to_bit(REQ_28) and (
	                       ( not k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and not k28_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and     k28_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k28_needs_attention) );

	k29_being_served <= to_bit(REQ_29) and (
	                       ( not k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and not bram_0_input_sel(1) and     bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and not bram_1_input_sel(1) and     bram_1_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and not bram_2_input_sel(1) and     bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and not bram_3_input_sel(1) and     bram_3_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and not bram_4_input_sel(1) and     bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and not bram_5_input_sel(1) and     bram_5_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and not bram_6_input_sel(1) and     bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and not bram_7_input_sel(1) and     bram_7_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and not bram_8_input_sel(1) and     bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and not bram_9_input_sel(1) and     bram_9_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and not bram_10_input_sel(1) and     bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and not bram_11_input_sel(1) and     bram_11_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and not bram_12_input_sel(1) and     bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and not bram_13_input_sel(1) and     bram_13_input_sel(0)) ) )
	                       or
	                       ( not k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and not bram_14_input_sel(1) and     bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and not bram_15_input_sel(1) and     bram_15_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and not bram_16_input_sel(1) and     bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and not bram_17_input_sel(1) and     bram_17_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and not bram_18_input_sel(1) and     bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and not bram_19_input_sel(1) and     bram_19_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and not bram_20_input_sel(1) and     bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and not bram_21_input_sel(1) and     bram_21_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and not bram_22_input_sel(1) and     bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and not bram_23_input_sel(1) and     bram_23_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and not bram_24_input_sel(1) and     bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and not bram_25_input_sel(1) and     bram_25_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and not bram_26_input_sel(1) and     bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and not bram_27_input_sel(1) and     bram_27_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and not k29_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and not bram_28_input_sel(1) and     bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and not bram_29_input_sel(1) and     bram_29_input_sel(0)) ) )
	                       or
	                       (     k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and     k29_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and not bram_30_input_sel(1) and     bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and not bram_31_input_sel(1) and     bram_31_input_sel(0)) ) )
	                       or
	                       (not k29_needs_attention) );

	k30_being_served <= to_bit(REQ_30) and (
	                       ( not k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_0_input_sel(4) and     bram_0_input_sel(3) and     bram_0_input_sel(2) and     bram_0_input_sel(1) and not bram_0_input_sel(0)) or
	                                                                             (     bram_1_input_sel(4) and     bram_1_input_sel(3) and     bram_1_input_sel(2) and     bram_1_input_sel(1) and not bram_1_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_2_input_sel(4) and     bram_2_input_sel(3) and     bram_2_input_sel(2) and     bram_2_input_sel(1) and not bram_2_input_sel(0)) or
	                                                                             (     bram_3_input_sel(4) and     bram_3_input_sel(3) and     bram_3_input_sel(2) and     bram_3_input_sel(1) and not bram_3_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_4_input_sel(4) and     bram_4_input_sel(3) and     bram_4_input_sel(2) and     bram_4_input_sel(1) and not bram_4_input_sel(0)) or
	                                                                             (     bram_5_input_sel(4) and     bram_5_input_sel(3) and     bram_5_input_sel(2) and     bram_5_input_sel(1) and not bram_5_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_6_input_sel(4) and     bram_6_input_sel(3) and     bram_6_input_sel(2) and     bram_6_input_sel(1) and not bram_6_input_sel(0)) or
	                                                                             (     bram_7_input_sel(4) and     bram_7_input_sel(3) and     bram_7_input_sel(2) and     bram_7_input_sel(1) and not bram_7_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_8_input_sel(4) and     bram_8_input_sel(3) and     bram_8_input_sel(2) and     bram_8_input_sel(1) and not bram_8_input_sel(0)) or
	                                                                             (     bram_9_input_sel(4) and     bram_9_input_sel(3) and     bram_9_input_sel(2) and     bram_9_input_sel(1) and not bram_9_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_10_input_sel(4) and     bram_10_input_sel(3) and     bram_10_input_sel(2) and     bram_10_input_sel(1) and not bram_10_input_sel(0)) or
	                                                                             (     bram_11_input_sel(4) and     bram_11_input_sel(3) and     bram_11_input_sel(2) and     bram_11_input_sel(1) and not bram_11_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_12_input_sel(4) and     bram_12_input_sel(3) and     bram_12_input_sel(2) and     bram_12_input_sel(1) and not bram_12_input_sel(0)) or
	                                                                             (     bram_13_input_sel(4) and     bram_13_input_sel(3) and     bram_13_input_sel(2) and     bram_13_input_sel(1) and not bram_13_input_sel(0)) ) )
	                       or
	                       ( not k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_14_input_sel(4) and     bram_14_input_sel(3) and     bram_14_input_sel(2) and     bram_14_input_sel(1) and not bram_14_input_sel(0)) or
	                                                                             (     bram_15_input_sel(4) and     bram_15_input_sel(3) and     bram_15_input_sel(2) and     bram_15_input_sel(1) and not bram_15_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_16_input_sel(4) and     bram_16_input_sel(3) and     bram_16_input_sel(2) and     bram_16_input_sel(1) and not bram_16_input_sel(0)) or
	                                                                             (     bram_17_input_sel(4) and     bram_17_input_sel(3) and     bram_17_input_sel(2) and     bram_17_input_sel(1) and not bram_17_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_18_input_sel(4) and     bram_18_input_sel(3) and     bram_18_input_sel(2) and     bram_18_input_sel(1) and not bram_18_input_sel(0)) or
	                                                                             (     bram_19_input_sel(4) and     bram_19_input_sel(3) and     bram_19_input_sel(2) and     bram_19_input_sel(1) and not bram_19_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_20_input_sel(4) and     bram_20_input_sel(3) and     bram_20_input_sel(2) and     bram_20_input_sel(1) and not bram_20_input_sel(0)) or
	                                                                             (     bram_21_input_sel(4) and     bram_21_input_sel(3) and     bram_21_input_sel(2) and     bram_21_input_sel(1) and not bram_21_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_22_input_sel(4) and     bram_22_input_sel(3) and     bram_22_input_sel(2) and     bram_22_input_sel(1) and not bram_22_input_sel(0)) or
	                                                                             (     bram_23_input_sel(4) and     bram_23_input_sel(3) and     bram_23_input_sel(2) and     bram_23_input_sel(1) and not bram_23_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_24_input_sel(4) and     bram_24_input_sel(3) and     bram_24_input_sel(2) and     bram_24_input_sel(1) and not bram_24_input_sel(0)) or
	                                                                             (     bram_25_input_sel(4) and     bram_25_input_sel(3) and     bram_25_input_sel(2) and     bram_25_input_sel(1) and not bram_25_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_26_input_sel(4) and     bram_26_input_sel(3) and     bram_26_input_sel(2) and     bram_26_input_sel(1) and not bram_26_input_sel(0)) or
	                                                                             (     bram_27_input_sel(4) and     bram_27_input_sel(3) and     bram_27_input_sel(2) and     bram_27_input_sel(1) and not bram_27_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and not k30_output_sel(0) and ( (     bram_28_input_sel(4) and     bram_28_input_sel(3) and     bram_28_input_sel(2) and     bram_28_input_sel(1) and not bram_28_input_sel(0)) or
	                                                                             (     bram_29_input_sel(4) and     bram_29_input_sel(3) and     bram_29_input_sel(2) and     bram_29_input_sel(1) and not bram_29_input_sel(0)) ) )
	                       or
	                       (     k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and     k30_output_sel(0) and ( (     bram_30_input_sel(4) and     bram_30_input_sel(3) and     bram_30_input_sel(2) and     bram_30_input_sel(1) and not bram_30_input_sel(0)) or
	                                                                             (     bram_31_input_sel(4) and     bram_31_input_sel(3) and     bram_31_input_sel(2) and     bram_31_input_sel(1) and not bram_31_input_sel(0)) ) )
	                       or
	                       (not k30_needs_attention) );

	k31_being_served <= to_bit(REQ_31);


	k0_output_sel(4 downto 1) <= to_bitvector(ADDR_0(12 downto 9));
	k1_output_sel(4 downto 1) <= to_bitvector(ADDR_1(12 downto 9));
	k2_output_sel(4 downto 1) <= to_bitvector(ADDR_2(12 downto 9));
	k3_output_sel(4 downto 1) <= to_bitvector(ADDR_3(12 downto 9));
	k4_output_sel(4 downto 1) <= to_bitvector(ADDR_4(12 downto 9));
	k5_output_sel(4 downto 1) <= to_bitvector(ADDR_5(12 downto 9));
	k6_output_sel(4 downto 1) <= to_bitvector(ADDR_6(12 downto 9));
	k7_output_sel(4 downto 1) <= to_bitvector(ADDR_7(12 downto 9));
	k8_output_sel(4 downto 1) <= to_bitvector(ADDR_8(12 downto 9));
	k9_output_sel(4 downto 1) <= to_bitvector(ADDR_9(12 downto 9));
	k10_output_sel(4 downto 1) <= to_bitvector(ADDR_10(12 downto 9));
	k11_output_sel(4 downto 1) <= to_bitvector(ADDR_11(12 downto 9));
	k12_output_sel(4 downto 1) <= to_bitvector(ADDR_12(12 downto 9));
	k13_output_sel(4 downto 1) <= to_bitvector(ADDR_13(12 downto 9));
	k14_output_sel(4 downto 1) <= to_bitvector(ADDR_14(12 downto 9));
	k15_output_sel(4 downto 1) <= to_bitvector(ADDR_15(12 downto 9));
	k16_output_sel(4 downto 1) <= to_bitvector(ADDR_16(12 downto 9));
	k17_output_sel(4 downto 1) <= to_bitvector(ADDR_17(12 downto 9));
	k18_output_sel(4 downto 1) <= to_bitvector(ADDR_18(12 downto 9));
	k19_output_sel(4 downto 1) <= to_bitvector(ADDR_19(12 downto 9));
	k20_output_sel(4 downto 1) <= to_bitvector(ADDR_20(12 downto 9));
	k21_output_sel(4 downto 1) <= to_bitvector(ADDR_21(12 downto 9));
	k22_output_sel(4 downto 1) <= to_bitvector(ADDR_22(12 downto 9));
	k23_output_sel(4 downto 1) <= to_bitvector(ADDR_23(12 downto 9));
	k24_output_sel(4 downto 1) <= to_bitvector(ADDR_24(12 downto 9));
	k25_output_sel(4 downto 1) <= to_bitvector(ADDR_25(12 downto 9));
	k26_output_sel(4 downto 1) <= to_bitvector(ADDR_26(12 downto 9));
	k27_output_sel(4 downto 1) <= to_bitvector(ADDR_27(12 downto 9));
	k28_output_sel(4 downto 1) <= to_bitvector(ADDR_28(12 downto 9));
	k29_output_sel(4 downto 1) <= to_bitvector(ADDR_29(12 downto 9));
	k30_output_sel(4 downto 1) <= to_bitvector(ADDR_30(12 downto 9));
	k31_output_sel(4 downto 1) <= to_bitvector(ADDR_31(12 downto 9));


	k0_output_sel(0) <= ( not k0_output_sel(4) and not k0_output_sel(3) and not k0_output_sel(2) and not k0_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and not k0_output_sel(3) and not k0_output_sel(2) and     k0_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and not k0_output_sel(3) and     k0_output_sel(2) and not k0_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and not k0_output_sel(3) and     k0_output_sel(2) and     k0_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and     k0_output_sel(3) and not k0_output_sel(2) and not k0_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and     k0_output_sel(3) and not k0_output_sel(2) and     k0_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and     k0_output_sel(3) and     k0_output_sel(2) and not k0_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k0_output_sel(4) and     k0_output_sel(3) and     k0_output_sel(2) and     k0_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and not k0_output_sel(3) and not k0_output_sel(2) and not k0_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and not k0_output_sel(3) and not k0_output_sel(2) and     k0_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and not k0_output_sel(3) and     k0_output_sel(2) and not k0_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and not k0_output_sel(3) and     k0_output_sel(2) and     k0_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and     k0_output_sel(3) and not k0_output_sel(2) and not k0_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and     k0_output_sel(3) and not k0_output_sel(2) and     k0_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and     k0_output_sel(3) and     k0_output_sel(2) and not k0_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k0_output_sel(4) and     k0_output_sel(3) and     k0_output_sel(2) and     k0_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k1_output_sel(0) <= ( not k1_output_sel(4) and not k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and not k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and not k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and not k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and     k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and     k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and     k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k1_output_sel(4) and     k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and not k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and not k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and not k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and not k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and     k1_output_sel(3) and not k1_output_sel(2) and not k1_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and     k1_output_sel(3) and not k1_output_sel(2) and     k1_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and     k1_output_sel(3) and     k1_output_sel(2) and not k1_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k1_output_sel(4) and     k1_output_sel(3) and     k1_output_sel(2) and     k1_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k2_output_sel(0) <= ( not k2_output_sel(4) and not k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and not k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and not k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and not k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and     k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and     k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and     k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k2_output_sel(4) and     k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and not k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and not k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and not k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and not k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and     k2_output_sel(3) and not k2_output_sel(2) and not k2_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and     k2_output_sel(3) and not k2_output_sel(2) and     k2_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and     k2_output_sel(3) and     k2_output_sel(2) and not k2_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k2_output_sel(4) and     k2_output_sel(3) and     k2_output_sel(2) and     k2_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k3_output_sel(0) <= ( not k3_output_sel(4) and not k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and not k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and not k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and not k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and     k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and     k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and     k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k3_output_sel(4) and     k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and not k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and not k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and not k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and not k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and     k3_output_sel(3) and not k3_output_sel(2) and not k3_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and     k3_output_sel(3) and not k3_output_sel(2) and     k3_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and     k3_output_sel(3) and     k3_output_sel(2) and not k3_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k3_output_sel(4) and     k3_output_sel(3) and     k3_output_sel(2) and     k3_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k4_output_sel(0) <= ( not k4_output_sel(4) and not k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and not k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and not k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and not k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and     k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and     k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and     k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k4_output_sel(4) and     k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and not k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and not k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and not k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and not k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and     k4_output_sel(3) and not k4_output_sel(2) and not k4_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and     k4_output_sel(3) and not k4_output_sel(2) and     k4_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and     k4_output_sel(3) and     k4_output_sel(2) and not k4_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k4_output_sel(4) and     k4_output_sel(3) and     k4_output_sel(2) and     k4_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k5_output_sel(0) <= ( not k5_output_sel(4) and not k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and not k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and not k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and not k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and     k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and     k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and     k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k5_output_sel(4) and     k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and not k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and not k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and not k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and not k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and     k5_output_sel(3) and not k5_output_sel(2) and not k5_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and     k5_output_sel(3) and not k5_output_sel(2) and     k5_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and     k5_output_sel(3) and     k5_output_sel(2) and not k5_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k5_output_sel(4) and     k5_output_sel(3) and     k5_output_sel(2) and     k5_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k6_output_sel(0) <= ( not k6_output_sel(4) and not k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and not k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and not k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and not k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and     k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and     k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and     k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k6_output_sel(4) and     k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and not k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and not k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and not k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and not k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and     k6_output_sel(3) and not k6_output_sel(2) and not k6_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and     k6_output_sel(3) and not k6_output_sel(2) and     k6_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and     k6_output_sel(3) and     k6_output_sel(2) and not k6_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k6_output_sel(4) and     k6_output_sel(3) and     k6_output_sel(2) and     k6_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k7_output_sel(0) <= ( not k7_output_sel(4) and not k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and not k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and not k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and not k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and     k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and     k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and     k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k7_output_sel(4) and     k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and not k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and not k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and not k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and not k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and     k7_output_sel(3) and not k7_output_sel(2) and not k7_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and     k7_output_sel(3) and not k7_output_sel(2) and     k7_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and     k7_output_sel(3) and     k7_output_sel(2) and not k7_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k7_output_sel(4) and     k7_output_sel(3) and     k7_output_sel(2) and     k7_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k8_output_sel(0) <= ( not k8_output_sel(4) and not k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and not k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and not k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and not k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and     k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and     k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and     k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k8_output_sel(4) and     k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and not k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and not k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and not k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and not k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and     k8_output_sel(3) and not k8_output_sel(2) and not k8_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and     k8_output_sel(3) and not k8_output_sel(2) and     k8_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and     k8_output_sel(3) and     k8_output_sel(2) and not k8_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k8_output_sel(4) and     k8_output_sel(3) and     k8_output_sel(2) and     k8_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k9_output_sel(0) <= ( not k9_output_sel(4) and not k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and not k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and not k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and not k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and     k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and     k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and     k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k9_output_sel(4) and     k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and not k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and not k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and not k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and not k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and     k9_output_sel(3) and not k9_output_sel(2) and not k9_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and     k9_output_sel(3) and not k9_output_sel(2) and     k9_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and     k9_output_sel(3) and     k9_output_sel(2) and not k9_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k9_output_sel(4) and     k9_output_sel(3) and     k9_output_sel(2) and     k9_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k10_output_sel(0) <= ( not k10_output_sel(4) and not k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and not k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and not k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and not k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and     k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and     k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and     k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k10_output_sel(4) and     k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and not k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and not k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and not k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and not k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and     k10_output_sel(3) and not k10_output_sel(2) and not k10_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and     k10_output_sel(3) and not k10_output_sel(2) and     k10_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and     k10_output_sel(3) and     k10_output_sel(2) and not k10_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k10_output_sel(4) and     k10_output_sel(3) and     k10_output_sel(2) and     k10_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k11_output_sel(0) <= ( not k11_output_sel(4) and not k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and not k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and not k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and not k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and     k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and     k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and     k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k11_output_sel(4) and     k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and not k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and not k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and not k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and not k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and     k11_output_sel(3) and not k11_output_sel(2) and not k11_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and     k11_output_sel(3) and not k11_output_sel(2) and     k11_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and     k11_output_sel(3) and     k11_output_sel(2) and not k11_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k11_output_sel(4) and     k11_output_sel(3) and     k11_output_sel(2) and     k11_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k12_output_sel(0) <= ( not k12_output_sel(4) and not k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and not k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and not k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and not k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and     k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and     k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and     k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k12_output_sel(4) and     k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and not k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and not k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and not k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and not k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and     k12_output_sel(3) and not k12_output_sel(2) and not k12_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and     k12_output_sel(3) and not k12_output_sel(2) and     k12_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and     k12_output_sel(3) and     k12_output_sel(2) and not k12_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k12_output_sel(4) and     k12_output_sel(3) and     k12_output_sel(2) and     k12_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k13_output_sel(0) <= ( not k13_output_sel(4) and not k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and not k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and not k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and not k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and     k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and     k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and     k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k13_output_sel(4) and     k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and not k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and not k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and not k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and not k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and     k13_output_sel(3) and not k13_output_sel(2) and not k13_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and     k13_output_sel(3) and not k13_output_sel(2) and     k13_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and     k13_output_sel(3) and     k13_output_sel(2) and not k13_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k13_output_sel(4) and     k13_output_sel(3) and     k13_output_sel(2) and     k13_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k14_output_sel(0) <= ( not k14_output_sel(4) and not k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and not k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and not k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and not k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and     k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and     k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and     k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k14_output_sel(4) and     k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and not k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and not k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and not k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and not k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and     k14_output_sel(3) and not k14_output_sel(2) and not k14_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and     k14_output_sel(3) and not k14_output_sel(2) and     k14_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and     k14_output_sel(3) and     k14_output_sel(2) and not k14_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k14_output_sel(4) and     k14_output_sel(3) and     k14_output_sel(2) and     k14_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k15_output_sel(0) <= ( not k15_output_sel(4) and not k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and ( not bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and not k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and ( not bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and not k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and ( not bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and not k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and ( not bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and     k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and ( not bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and     k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and ( not bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and     k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and ( not bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k15_output_sel(4) and     k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and ( not bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and not k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and ( not bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and not k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and ( not bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and not k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and ( not bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and not k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and ( not bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and     k15_output_sel(3) and not k15_output_sel(2) and not k15_output_sel(1) and ( not bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and     k15_output_sel(3) and not k15_output_sel(2) and     k15_output_sel(1) and ( not bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and     k15_output_sel(3) and     k15_output_sel(2) and not k15_output_sel(1) and ( not bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k15_output_sel(4) and     k15_output_sel(3) and     k15_output_sel(2) and     k15_output_sel(1) and ( not bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k16_output_sel(0) <= ( not k16_output_sel(4) and not k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and not k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and not k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and not k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and     k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and     k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and     k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k16_output_sel(4) and     k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and not k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and not k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and not k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and not k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and     k16_output_sel(3) and not k16_output_sel(2) and not k16_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and     k16_output_sel(3) and not k16_output_sel(2) and     k16_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and     k16_output_sel(3) and     k16_output_sel(2) and not k16_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k16_output_sel(4) and     k16_output_sel(3) and     k16_output_sel(2) and     k16_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k17_output_sel(0) <= ( not k17_output_sel(4) and not k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and not k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and not k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and not k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and     k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and     k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and     k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k17_output_sel(4) and     k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and not k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and not k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and not k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and not k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and     k17_output_sel(3) and not k17_output_sel(2) and not k17_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and     k17_output_sel(3) and not k17_output_sel(2) and     k17_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and     k17_output_sel(3) and     k17_output_sel(2) and not k17_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k17_output_sel(4) and     k17_output_sel(3) and     k17_output_sel(2) and     k17_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k18_output_sel(0) <= ( not k18_output_sel(4) and not k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and not k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and not k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and not k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and     k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and     k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and     k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k18_output_sel(4) and     k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and not k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and not k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and not k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and not k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and     k18_output_sel(3) and not k18_output_sel(2) and not k18_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and     k18_output_sel(3) and not k18_output_sel(2) and     k18_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and     k18_output_sel(3) and     k18_output_sel(2) and not k18_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k18_output_sel(4) and     k18_output_sel(3) and     k18_output_sel(2) and     k18_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k19_output_sel(0) <= ( not k19_output_sel(4) and not k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and not k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and not k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and not k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and     k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and     k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and     k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k19_output_sel(4) and     k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and not k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and not k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and not k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and not k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and     k19_output_sel(3) and not k19_output_sel(2) and not k19_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and     k19_output_sel(3) and not k19_output_sel(2) and     k19_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and     k19_output_sel(3) and     k19_output_sel(2) and not k19_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k19_output_sel(4) and     k19_output_sel(3) and     k19_output_sel(2) and     k19_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k20_output_sel(0) <= ( not k20_output_sel(4) and not k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and not k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and not k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and not k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and     k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and     k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and     k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k20_output_sel(4) and     k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and not k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and not k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and not k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and not k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and     k20_output_sel(3) and not k20_output_sel(2) and not k20_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and     k20_output_sel(3) and not k20_output_sel(2) and     k20_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and     k20_output_sel(3) and     k20_output_sel(2) and not k20_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k20_output_sel(4) and     k20_output_sel(3) and     k20_output_sel(2) and     k20_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k21_output_sel(0) <= ( not k21_output_sel(4) and not k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and not k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and not k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and not k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and     k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and     k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and     k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k21_output_sel(4) and     k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and not k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and not k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and not k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and not k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and     k21_output_sel(3) and not k21_output_sel(2) and not k21_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and     k21_output_sel(3) and not k21_output_sel(2) and     k21_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and     k21_output_sel(3) and     k21_output_sel(2) and not k21_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k21_output_sel(4) and     k21_output_sel(3) and     k21_output_sel(2) and     k21_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k22_output_sel(0) <= ( not k22_output_sel(4) and not k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and not k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and not k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and not k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and     k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and     k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and     k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k22_output_sel(4) and     k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and not k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and not k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and not k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and not k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and     k22_output_sel(3) and not k22_output_sel(2) and not k22_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and     k22_output_sel(3) and not k22_output_sel(2) and     k22_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and     k22_output_sel(3) and     k22_output_sel(2) and not k22_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k22_output_sel(4) and     k22_output_sel(3) and     k22_output_sel(2) and     k22_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k23_output_sel(0) <= ( not k23_output_sel(4) and not k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                          not bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and not k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                          not bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and not k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                          not bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and not k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                          not bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and     k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                          not bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and     k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                          not bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and     k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                          not bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k23_output_sel(4) and     k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                          not bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and not k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                          not bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and not k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                          not bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and not k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                          not bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and not k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                          not bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and     k23_output_sel(3) and not k23_output_sel(2) and not k23_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                          not bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and     k23_output_sel(3) and not k23_output_sel(2) and     k23_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                          not bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and     k23_output_sel(3) and     k23_output_sel(2) and not k23_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                          not bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k23_output_sel(4) and     k23_output_sel(3) and     k23_output_sel(2) and     k23_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                          not bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k24_output_sel(0) <= ( not k24_output_sel(4) and not k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and not k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and not k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and not k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and     k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and     k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and     k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k24_output_sel(4) and     k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and not k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and not k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and not k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and not k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and     k24_output_sel(3) and not k24_output_sel(2) and not k24_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and     k24_output_sel(3) and not k24_output_sel(2) and     k24_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and     k24_output_sel(3) and     k24_output_sel(2) and not k24_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k24_output_sel(4) and     k24_output_sel(3) and     k24_output_sel(2) and     k24_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k25_output_sel(0) <= ( not k25_output_sel(4) and not k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and not k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and not k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and not k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and     k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and     k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and     k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k25_output_sel(4) and     k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and not k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and not k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and not k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and not k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and     k25_output_sel(3) and not k25_output_sel(2) and not k25_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and     k25_output_sel(3) and not k25_output_sel(2) and     k25_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and     k25_output_sel(3) and     k25_output_sel(2) and not k25_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k25_output_sel(4) and     k25_output_sel(3) and     k25_output_sel(2) and     k25_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k26_output_sel(0) <= ( not k26_output_sel(4) and not k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and not k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and not k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and not k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and     k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and     k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and     k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k26_output_sel(4) and     k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and not k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and not k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and not k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and not k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and     k26_output_sel(3) and not k26_output_sel(2) and not k26_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and     k26_output_sel(3) and not k26_output_sel(2) and     k26_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and     k26_output_sel(3) and     k26_output_sel(2) and not k26_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k26_output_sel(4) and     k26_output_sel(3) and     k26_output_sel(2) and     k26_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k27_output_sel(0) <= ( not k27_output_sel(4) and not k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                          not bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and not k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                          not bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and not k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                          not bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and not k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                          not bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and     k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                          not bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and     k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                          not bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and     k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                          not bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k27_output_sel(4) and     k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                          not bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and not k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                          not bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and not k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                          not bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and not k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                          not bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and not k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                          not bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and     k27_output_sel(3) and not k27_output_sel(2) and not k27_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                          not bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and     k27_output_sel(3) and not k27_output_sel(2) and     k27_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                          not bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and     k27_output_sel(3) and     k27_output_sel(2) and not k27_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                          not bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k27_output_sel(4) and     k27_output_sel(3) and     k27_output_sel(2) and     k27_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                          not bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k28_output_sel(0) <= ( not k28_output_sel(4) and not k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and not k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and not k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and not k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and     k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and     k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and     k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k28_output_sel(4) and     k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and not k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and not k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and not k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and not k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and     k28_output_sel(3) and not k28_output_sel(2) and not k28_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and     k28_output_sel(3) and not k28_output_sel(2) and     k28_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and     k28_output_sel(3) and     k28_output_sel(2) and not k28_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k28_output_sel(4) and     k28_output_sel(3) and     k28_output_sel(2) and     k28_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k29_output_sel(0) <= ( not k29_output_sel(4) and not k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                          not bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and not k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                          not bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and not k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                          not bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and not k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                          not bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and     k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                          not bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and     k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                          not bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and     k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                          not bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k29_output_sel(4) and     k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                          not bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and not k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                          not bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and not k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                          not bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and not k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                          not bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and not k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                          not bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and     k29_output_sel(3) and not k29_output_sel(2) and not k29_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                          not bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and     k29_output_sel(3) and not k29_output_sel(2) and     k29_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                          not bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and     k29_output_sel(3) and     k29_output_sel(2) and not k29_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                          not bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k29_output_sel(4) and     k29_output_sel(3) and     k29_output_sel(2) and     k29_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                          not bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );

	k30_output_sel(0) <= ( not k30_output_sel(4) and not k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                          not bram_1_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and not k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                          not bram_3_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and not k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                          not bram_5_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and not k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                          not bram_7_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and     k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                          not bram_9_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and     k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                          not bram_11_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and     k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                          not bram_13_input_sel(0)) )
	                    or
	                    ( not k30_output_sel(4) and     k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                          not bram_15_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and not k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                          not bram_17_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and not k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                          not bram_19_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and not k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                          not bram_21_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and not k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                          not bram_23_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and     k30_output_sel(3) and not k30_output_sel(2) and not k30_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                          not bram_25_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and     k30_output_sel(3) and not k30_output_sel(2) and     k30_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                          not bram_27_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and     k30_output_sel(3) and     k30_output_sel(2) and not k30_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                          not bram_29_input_sel(0)) )
	                    or
	                    (     k30_output_sel(4) and     k30_output_sel(3) and     k30_output_sel(2) and     k30_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                          not bram_31_input_sel(0)) );

	k31_output_sel(0) <= ( not k31_output_sel(4) and not k31_output_sel(3) and not k31_output_sel(2) and not k31_output_sel(1) and (     bram_1_input_sel(4) and
	                                                                              bram_1_input_sel(3) and
	                                                                              bram_1_input_sel(2) and
	                                                                              bram_1_input_sel(1) and
	                                                                              bram_1_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and not k31_output_sel(3) and not k31_output_sel(2) and     k31_output_sel(1) and (     bram_3_input_sel(4) and
	                                                                              bram_3_input_sel(3) and
	                                                                              bram_3_input_sel(2) and
	                                                                              bram_3_input_sel(1) and
	                                                                              bram_3_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and not k31_output_sel(3) and     k31_output_sel(2) and not k31_output_sel(1) and (     bram_5_input_sel(4) and
	                                                                              bram_5_input_sel(3) and
	                                                                              bram_5_input_sel(2) and
	                                                                              bram_5_input_sel(1) and
	                                                                              bram_5_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and not k31_output_sel(3) and     k31_output_sel(2) and     k31_output_sel(1) and (     bram_7_input_sel(4) and
	                                                                              bram_7_input_sel(3) and
	                                                                              bram_7_input_sel(2) and
	                                                                              bram_7_input_sel(1) and
	                                                                              bram_7_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and     k31_output_sel(3) and not k31_output_sel(2) and not k31_output_sel(1) and (     bram_9_input_sel(4) and
	                                                                              bram_9_input_sel(3) and
	                                                                              bram_9_input_sel(2) and
	                                                                              bram_9_input_sel(1) and
	                                                                              bram_9_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and     k31_output_sel(3) and not k31_output_sel(2) and     k31_output_sel(1) and (     bram_11_input_sel(4) and
	                                                                              bram_11_input_sel(3) and
	                                                                              bram_11_input_sel(2) and
	                                                                              bram_11_input_sel(1) and
	                                                                              bram_11_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and     k31_output_sel(3) and     k31_output_sel(2) and not k31_output_sel(1) and (     bram_13_input_sel(4) and
	                                                                              bram_13_input_sel(3) and
	                                                                              bram_13_input_sel(2) and
	                                                                              bram_13_input_sel(1) and
	                                                                              bram_13_input_sel(0)) )
	                    or
	                    ( not k31_output_sel(4) and     k31_output_sel(3) and     k31_output_sel(2) and     k31_output_sel(1) and (     bram_15_input_sel(4) and
	                                                                              bram_15_input_sel(3) and
	                                                                              bram_15_input_sel(2) and
	                                                                              bram_15_input_sel(1) and
	                                                                              bram_15_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and not k31_output_sel(3) and not k31_output_sel(2) and not k31_output_sel(1) and (     bram_17_input_sel(4) and
	                                                                              bram_17_input_sel(3) and
	                                                                              bram_17_input_sel(2) and
	                                                                              bram_17_input_sel(1) and
	                                                                              bram_17_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and not k31_output_sel(3) and not k31_output_sel(2) and     k31_output_sel(1) and (     bram_19_input_sel(4) and
	                                                                              bram_19_input_sel(3) and
	                                                                              bram_19_input_sel(2) and
	                                                                              bram_19_input_sel(1) and
	                                                                              bram_19_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and not k31_output_sel(3) and     k31_output_sel(2) and not k31_output_sel(1) and (     bram_21_input_sel(4) and
	                                                                              bram_21_input_sel(3) and
	                                                                              bram_21_input_sel(2) and
	                                                                              bram_21_input_sel(1) and
	                                                                              bram_21_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and not k31_output_sel(3) and     k31_output_sel(2) and     k31_output_sel(1) and (     bram_23_input_sel(4) and
	                                                                              bram_23_input_sel(3) and
	                                                                              bram_23_input_sel(2) and
	                                                                              bram_23_input_sel(1) and
	                                                                              bram_23_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and     k31_output_sel(3) and not k31_output_sel(2) and not k31_output_sel(1) and (     bram_25_input_sel(4) and
	                                                                              bram_25_input_sel(3) and
	                                                                              bram_25_input_sel(2) and
	                                                                              bram_25_input_sel(1) and
	                                                                              bram_25_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and     k31_output_sel(3) and not k31_output_sel(2) and     k31_output_sel(1) and (     bram_27_input_sel(4) and
	                                                                              bram_27_input_sel(3) and
	                                                                              bram_27_input_sel(2) and
	                                                                              bram_27_input_sel(1) and
	                                                                              bram_27_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and     k31_output_sel(3) and     k31_output_sel(2) and not k31_output_sel(1) and (     bram_29_input_sel(4) and
	                                                                              bram_29_input_sel(3) and
	                                                                              bram_29_input_sel(2) and
	                                                                              bram_29_input_sel(1) and
	                                                                              bram_29_input_sel(0)) )
	                    or
	                    (     k31_output_sel(4) and     k31_output_sel(3) and     k31_output_sel(2) and     k31_output_sel(1) and (     bram_31_input_sel(4) and
	                                                                              bram_31_input_sel(3) and
	                                                                              bram_31_input_sel(2) and
	                                                                              bram_31_input_sel(1) and
	                                                                              bram_31_input_sel(0)) );


	input_controller_0 : block begin
		with bram_0_input_sel select
			bram_di(1 * 32 - 1 downto 0 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_0_input_sel select
			bram_addr(1 * 9 - 1 downto 0 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_0_input_sel select
			bram_we(1 * 4 - 1 downto 0 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_0;

	input_controller_1 : block begin
		with bram_1_input_sel select
			bram_di(2 * 32 - 1 downto 1 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_1_input_sel select
			bram_addr(2 * 9 - 1 downto 1 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_1_input_sel select
			bram_we(2 * 4 - 1 downto 1 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_1;

	input_controller_2 : block begin
		with bram_2_input_sel select
			bram_di(3 * 32 - 1 downto 2 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_2_input_sel select
			bram_addr(3 * 9 - 1 downto 2 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_2_input_sel select
			bram_we(3 * 4 - 1 downto 2 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_2;

	input_controller_3 : block begin
		with bram_3_input_sel select
			bram_di(4 * 32 - 1 downto 3 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_3_input_sel select
			bram_addr(4 * 9 - 1 downto 3 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_3_input_sel select
			bram_we(4 * 4 - 1 downto 3 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_3;

	input_controller_4 : block begin
		with bram_4_input_sel select
			bram_di(5 * 32 - 1 downto 4 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_4_input_sel select
			bram_addr(5 * 9 - 1 downto 4 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_4_input_sel select
			bram_we(5 * 4 - 1 downto 4 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_4;

	input_controller_5 : block begin
		with bram_5_input_sel select
			bram_di(6 * 32 - 1 downto 5 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_5_input_sel select
			bram_addr(6 * 9 - 1 downto 5 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_5_input_sel select
			bram_we(6 * 4 - 1 downto 5 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_5;

	input_controller_6 : block begin
		with bram_6_input_sel select
			bram_di(7 * 32 - 1 downto 6 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_6_input_sel select
			bram_addr(7 * 9 - 1 downto 6 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_6_input_sel select
			bram_we(7 * 4 - 1 downto 6 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_6;

	input_controller_7 : block begin
		with bram_7_input_sel select
			bram_di(8 * 32 - 1 downto 7 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_7_input_sel select
			bram_addr(8 * 9 - 1 downto 7 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_7_input_sel select
			bram_we(8 * 4 - 1 downto 7 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_7;

	input_controller_8 : block begin
		with bram_8_input_sel select
			bram_di(9 * 32 - 1 downto 8 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_8_input_sel select
			bram_addr(9 * 9 - 1 downto 8 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_8_input_sel select
			bram_we(9 * 4 - 1 downto 8 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_8;

	input_controller_9 : block begin
		with bram_9_input_sel select
			bram_di(10 * 32 - 1 downto 9 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_9_input_sel select
			bram_addr(10 * 9 - 1 downto 9 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_9_input_sel select
			bram_we(10 * 4 - 1 downto 9 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_9;

	input_controller_10 : block begin
		with bram_10_input_sel select
			bram_di(11 * 32 - 1 downto 10 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_10_input_sel select
			bram_addr(11 * 9 - 1 downto 10 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_10_input_sel select
			bram_we(11 * 4 - 1 downto 10 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_10;

	input_controller_11 : block begin
		with bram_11_input_sel select
			bram_di(12 * 32 - 1 downto 11 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_11_input_sel select
			bram_addr(12 * 9 - 1 downto 11 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_11_input_sel select
			bram_we(12 * 4 - 1 downto 11 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_11;

	input_controller_12 : block begin
		with bram_12_input_sel select
			bram_di(13 * 32 - 1 downto 12 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_12_input_sel select
			bram_addr(13 * 9 - 1 downto 12 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_12_input_sel select
			bram_we(13 * 4 - 1 downto 12 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_12;

	input_controller_13 : block begin
		with bram_13_input_sel select
			bram_di(14 * 32 - 1 downto 13 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_13_input_sel select
			bram_addr(14 * 9 - 1 downto 13 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_13_input_sel select
			bram_we(14 * 4 - 1 downto 13 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_13;

	input_controller_14 : block begin
		with bram_14_input_sel select
			bram_di(15 * 32 - 1 downto 14 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_14_input_sel select
			bram_addr(15 * 9 - 1 downto 14 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_14_input_sel select
			bram_we(15 * 4 - 1 downto 14 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_14;

	input_controller_15 : block begin
		with bram_15_input_sel select
			bram_di(16 * 32 - 1 downto 15 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_15_input_sel select
			bram_addr(16 * 9 - 1 downto 15 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_15_input_sel select
			bram_we(16 * 4 - 1 downto 15 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_15;

	input_controller_16 : block begin
		with bram_16_input_sel select
			bram_di(17 * 32 - 1 downto 16 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_16_input_sel select
			bram_addr(17 * 9 - 1 downto 16 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_16_input_sel select
			bram_we(17 * 4 - 1 downto 16 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_16;

	input_controller_17 : block begin
		with bram_17_input_sel select
			bram_di(18 * 32 - 1 downto 17 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_17_input_sel select
			bram_addr(18 * 9 - 1 downto 17 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_17_input_sel select
			bram_we(18 * 4 - 1 downto 17 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_17;

	input_controller_18 : block begin
		with bram_18_input_sel select
			bram_di(19 * 32 - 1 downto 18 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_18_input_sel select
			bram_addr(19 * 9 - 1 downto 18 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_18_input_sel select
			bram_we(19 * 4 - 1 downto 18 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_18;

	input_controller_19 : block begin
		with bram_19_input_sel select
			bram_di(20 * 32 - 1 downto 19 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_19_input_sel select
			bram_addr(20 * 9 - 1 downto 19 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_19_input_sel select
			bram_we(20 * 4 - 1 downto 19 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_19;

	input_controller_20 : block begin
		with bram_20_input_sel select
			bram_di(21 * 32 - 1 downto 20 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_20_input_sel select
			bram_addr(21 * 9 - 1 downto 20 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_20_input_sel select
			bram_we(21 * 4 - 1 downto 20 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_20;

	input_controller_21 : block begin
		with bram_21_input_sel select
			bram_di(22 * 32 - 1 downto 21 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_21_input_sel select
			bram_addr(22 * 9 - 1 downto 21 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_21_input_sel select
			bram_we(22 * 4 - 1 downto 21 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_21;

	input_controller_22 : block begin
		with bram_22_input_sel select
			bram_di(23 * 32 - 1 downto 22 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_22_input_sel select
			bram_addr(23 * 9 - 1 downto 22 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_22_input_sel select
			bram_we(23 * 4 - 1 downto 22 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_22;

	input_controller_23 : block begin
		with bram_23_input_sel select
			bram_di(24 * 32 - 1 downto 23 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_23_input_sel select
			bram_addr(24 * 9 - 1 downto 23 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_23_input_sel select
			bram_we(24 * 4 - 1 downto 23 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_23;

	input_controller_24 : block begin
		with bram_24_input_sel select
			bram_di(25 * 32 - 1 downto 24 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_24_input_sel select
			bram_addr(25 * 9 - 1 downto 24 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_24_input_sel select
			bram_we(25 * 4 - 1 downto 24 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_24;

	input_controller_25 : block begin
		with bram_25_input_sel select
			bram_di(26 * 32 - 1 downto 25 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_25_input_sel select
			bram_addr(26 * 9 - 1 downto 25 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_25_input_sel select
			bram_we(26 * 4 - 1 downto 25 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_25;

	input_controller_26 : block begin
		with bram_26_input_sel select
			bram_di(27 * 32 - 1 downto 26 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_26_input_sel select
			bram_addr(27 * 9 - 1 downto 26 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_26_input_sel select
			bram_we(27 * 4 - 1 downto 26 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_26;

	input_controller_27 : block begin
		with bram_27_input_sel select
			bram_di(28 * 32 - 1 downto 27 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_27_input_sel select
			bram_addr(28 * 9 - 1 downto 27 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_27_input_sel select
			bram_we(28 * 4 - 1 downto 27 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_27;

	input_controller_28 : block begin
		with bram_28_input_sel select
			bram_di(29 * 32 - 1 downto 28 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_28_input_sel select
			bram_addr(29 * 9 - 1 downto 28 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_28_input_sel select
			bram_we(29 * 4 - 1 downto 28 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_28;

	input_controller_29 : block begin
		with bram_29_input_sel select
			bram_di(30 * 32 - 1 downto 29 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_29_input_sel select
			bram_addr(30 * 9 - 1 downto 29 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_29_input_sel select
			bram_we(30 * 4 - 1 downto 29 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_29;

	input_controller_30 : block begin
		with bram_30_input_sel select
			bram_di(31 * 32 - 1 downto 30 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_30_input_sel select
			bram_addr(31 * 9 - 1 downto 30 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_30_input_sel select
			bram_we(31 * 4 - 1 downto 30 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_30;

	input_controller_31 : block begin
		with bram_31_input_sel select
			bram_di(32 * 32 - 1 downto 31 * 32)    <=  DI(32 * 1 - 1 downto 32 * 0) when "00000",
			              DI(32 * 2 - 1 downto 32 * 1) when "00001",
			              DI(32 * 3 - 1 downto 32 * 2) when "00010",
			              DI(32 * 4 - 1 downto 32 * 3) when "00011",
			              DI(32 * 5 - 1 downto 32 * 4) when "00100",
			              DI(32 * 6 - 1 downto 32 * 5) when "00101",
			              DI(32 * 7 - 1 downto 32 * 6) when "00110",
			              DI(32 * 8 - 1 downto 32 * 7) when "00111",
			              DI(32 * 9 - 1 downto 32 * 8) when "01000",
			              DI(32 * 10 - 1 downto 32 * 9) when "01001",
			              DI(32 * 11 - 1 downto 32 * 10) when "01010",
			              DI(32 * 12 - 1 downto 32 * 11) when "01011",
			              DI(32 * 13 - 1 downto 32 * 12) when "01100",
			              DI(32 * 14 - 1 downto 32 * 13) when "01101",
			              DI(32 * 15 - 1 downto 32 * 14) when "01110",
			              DI(32 * 16 - 1 downto 32 * 15) when "01111",
			              DI(32 * 17 - 1 downto 32 * 16) when "10000",
			              DI(32 * 18 - 1 downto 32 * 17) when "10001",
			              DI(32 * 19 - 1 downto 32 * 18) when "10010",
			              DI(32 * 20 - 1 downto 32 * 19) when "10011",
			              DI(32 * 21 - 1 downto 32 * 20) when "10100",
			              DI(32 * 22 - 1 downto 32 * 21) when "10101",
			              DI(32 * 23 - 1 downto 32 * 22) when "10110",
			              DI(32 * 24 - 1 downto 32 * 23) when "10111",
			              DI(32 * 25 - 1 downto 32 * 24) when "11000",
			              DI(32 * 26 - 1 downto 32 * 25) when "11001",
			              DI(32 * 27 - 1 downto 32 * 26) when "11010",
			              DI(32 * 28 - 1 downto 32 * 27) when "11011",
			              DI(32 * 29 - 1 downto 32 * 28) when "11100",
			              DI(32 * 30 - 1 downto 32 * 29) when "11101",
			              DI(32 * 31 - 1 downto 32 * 30) when "11110",
			              DI(32 * 32 - 1 downto 32 * 31) when "11111";
		with bram_31_input_sel select
			bram_addr(32 * 9 - 1 downto 31 * 9)  <=  ADDR_0(8 downto 0) when "00000",
			              ADDR_1(8 downto 0) when "00001",
			              ADDR_2(8 downto 0) when "00010",
			              ADDR_3(8 downto 0) when "00011",
			              ADDR_4(8 downto 0) when "00100",
			              ADDR_5(8 downto 0) when "00101",
			              ADDR_6(8 downto 0) when "00110",
			              ADDR_7(8 downto 0) when "00111",
			              ADDR_8(8 downto 0) when "01000",
			              ADDR_9(8 downto 0) when "01001",
			              ADDR_10(8 downto 0) when "01010",
			              ADDR_11(8 downto 0) when "01011",
			              ADDR_12(8 downto 0) when "01100",
			              ADDR_13(8 downto 0) when "01101",
			              ADDR_14(8 downto 0) when "01110",
			              ADDR_15(8 downto 0) when "01111",
			              ADDR_16(8 downto 0) when "10000",
			              ADDR_17(8 downto 0) when "10001",
			              ADDR_18(8 downto 0) when "10010",
			              ADDR_19(8 downto 0) when "10011",
			              ADDR_20(8 downto 0) when "10100",
			              ADDR_21(8 downto 0) when "10101",
			              ADDR_22(8 downto 0) when "10110",
			              ADDR_23(8 downto 0) when "10111",
			              ADDR_24(8 downto 0) when "11000",
			              ADDR_25(8 downto 0) when "11001",
			              ADDR_26(8 downto 0) when "11010",
			              ADDR_27(8 downto 0) when "11011",
			              ADDR_28(8 downto 0) when "11100",
			              ADDR_29(8 downto 0) when "11101",
			              ADDR_30(8 downto 0) when "11110",
			              ADDR_31(8 downto 0) when "11111";
		with bram_31_input_sel select
			bram_we(32 * 4 - 1 downto 31 * 4)    <=  we_0_safe when "00000",
			              we_1_safe when "00001",
			              we_2_safe when "00010",
			              we_3_safe when "00011",
			              we_4_safe when "00100",
			              we_5_safe when "00101",
			              we_6_safe when "00110",
			              we_7_safe when "00111",
			              we_8_safe when "01000",
			              we_9_safe when "01001",
			              we_10_safe when "01010",
			              we_11_safe when "01011",
			              we_12_safe when "01100",
			              we_13_safe when "01101",
			              we_14_safe when "01110",
			              we_15_safe when "01111",
			              we_16_safe when "10000",
			              we_17_safe when "10001",
			              we_18_safe when "10010",
			              we_19_safe when "10011",
			              we_20_safe when "10100",
			              we_21_safe when "10101",
			              we_22_safe when "10110",
			              we_23_safe when "10111",
			              we_24_safe when "11000",
			              we_25_safe when "11001",
			              we_26_safe when "11010",
			              we_27_safe when "11011",
			              we_28_safe when "11100",
			              we_29_safe when "11101",
			              we_30_safe when "11110",
			              we_31_safe when "11111";
	end block input_controller_31;


	output_controller_0 : block begin
		with k0_output_sel select
			DO(32 * 1 - 1 downto 32 * 0) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_0;

	output_controller_1 : block begin
		with k1_output_sel select
			DO(32 * 2 - 1 downto 32 * 1) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_1;

	output_controller_2 : block begin
		with k2_output_sel select
			DO(32 * 3 - 1 downto 32 * 2) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_2;

	output_controller_3 : block begin
		with k3_output_sel select
			DO(32 * 4 - 1 downto 32 * 3) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_3;

	output_controller_4 : block begin
		with k4_output_sel select
			DO(32 * 5 - 1 downto 32 * 4) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_4;

	output_controller_5 : block begin
		with k5_output_sel select
			DO(32 * 6 - 1 downto 32 * 5) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_5;

	output_controller_6 : block begin
		with k6_output_sel select
			DO(32 * 7 - 1 downto 32 * 6) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_6;

	output_controller_7 : block begin
		with k7_output_sel select
			DO(32 * 8 - 1 downto 32 * 7) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_7;

	output_controller_8 : block begin
		with k8_output_sel select
			DO(32 * 9 - 1 downto 32 * 8) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_8;

	output_controller_9 : block begin
		with k9_output_sel select
			DO(32 * 10 - 1 downto 32 * 9) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_9;

	output_controller_10 : block begin
		with k10_output_sel select
			DO(32 * 11 - 1 downto 32 * 10) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_10;

	output_controller_11 : block begin
		with k11_output_sel select
			DO(32 * 12 - 1 downto 32 * 11) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_11;

	output_controller_12 : block begin
		with k12_output_sel select
			DO(32 * 13 - 1 downto 32 * 12) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_12;

	output_controller_13 : block begin
		with k13_output_sel select
			DO(32 * 14 - 1 downto 32 * 13) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_13;

	output_controller_14 : block begin
		with k14_output_sel select
			DO(32 * 15 - 1 downto 32 * 14) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_14;

	output_controller_15 : block begin
		with k15_output_sel select
			DO(32 * 16 - 1 downto 32 * 15) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_15;

	output_controller_16 : block begin
		with k16_output_sel select
			DO(32 * 17 - 1 downto 32 * 16) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_16;

	output_controller_17 : block begin
		with k17_output_sel select
			DO(32 * 18 - 1 downto 32 * 17) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_17;

	output_controller_18 : block begin
		with k18_output_sel select
			DO(32 * 19 - 1 downto 32 * 18) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_18;

	output_controller_19 : block begin
		with k19_output_sel select
			DO(32 * 20 - 1 downto 32 * 19) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_19;

	output_controller_20 : block begin
		with k20_output_sel select
			DO(32 * 21 - 1 downto 32 * 20) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_20;

	output_controller_21 : block begin
		with k21_output_sel select
			DO(32 * 22 - 1 downto 32 * 21) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_21;

	output_controller_22 : block begin
		with k22_output_sel select
			DO(32 * 23 - 1 downto 32 * 22) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_22;

	output_controller_23 : block begin
		with k23_output_sel select
			DO(32 * 24 - 1 downto 32 * 23) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_23;

	output_controller_24 : block begin
		with k24_output_sel select
			DO(32 * 25 - 1 downto 32 * 24) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_24;

	output_controller_25 : block begin
		with k25_output_sel select
			DO(32 * 26 - 1 downto 32 * 25) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_25;

	output_controller_26 : block begin
		with k26_output_sel select
			DO(32 * 27 - 1 downto 32 * 26) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_26;

	output_controller_27 : block begin
		with k27_output_sel select
			DO(32 * 28 - 1 downto 32 * 27) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_27;

	output_controller_28 : block begin
		with k28_output_sel select
			DO(32 * 29 - 1 downto 32 * 28) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_28;

	output_controller_29 : block begin
		with k29_output_sel select
			DO(32 * 30 - 1 downto 32 * 29) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_29;

	output_controller_30 : block begin
		with k30_output_sel select
			DO(32 * 31 - 1 downto 32 * 30) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_30;

	output_controller_31 : block begin
		with k31_output_sel select
			DO(32 * 32 - 1 downto 32 * 31) <= bram_do(1 * 32 - 1 downto 0 * 32) when "00000",
			        bram_do(2 * 32 - 1 downto 1 * 32) when "00001",
			        bram_do(3 * 32 - 1 downto 2 * 32) when "00010",
			        bram_do(4 * 32 - 1 downto 3 * 32) when "00011",
			        bram_do(5 * 32 - 1 downto 4 * 32) when "00100",
			        bram_do(6 * 32 - 1 downto 5 * 32) when "00101",
			        bram_do(7 * 32 - 1 downto 6 * 32) when "00110",
			        bram_do(8 * 32 - 1 downto 7 * 32) when "00111",
			        bram_do(9 * 32 - 1 downto 8 * 32) when "01000",
			        bram_do(10 * 32 - 1 downto 9 * 32) when "01001",
			        bram_do(11 * 32 - 1 downto 10 * 32) when "01010",
			        bram_do(12 * 32 - 1 downto 11 * 32) when "01011",
			        bram_do(13 * 32 - 1 downto 12 * 32) when "01100",
			        bram_do(14 * 32 - 1 downto 13 * 32) when "01101",
			        bram_do(15 * 32 - 1 downto 14 * 32) when "01110",
			        bram_do(16 * 32 - 1 downto 15 * 32) when "01111",
			        bram_do(17 * 32 - 1 downto 16 * 32) when "10000",
			        bram_do(18 * 32 - 1 downto 17 * 32) when "10001",
			        bram_do(19 * 32 - 1 downto 18 * 32) when "10010",
			        bram_do(20 * 32 - 1 downto 19 * 32) when "10011",
			        bram_do(21 * 32 - 1 downto 20 * 32) when "10100",
			        bram_do(22 * 32 - 1 downto 21 * 32) when "10101",
			        bram_do(23 * 32 - 1 downto 22 * 32) when "10110",
			        bram_do(24 * 32 - 1 downto 23 * 32) when "10111",
			        bram_do(25 * 32 - 1 downto 24 * 32) when "11000",
			        bram_do(26 * 32 - 1 downto 25 * 32) when "11001",
			        bram_do(27 * 32 - 1 downto 26 * 32) when "11010",
			        bram_do(28 * 32 - 1 downto 27 * 32) when "11011",
			        bram_do(29 * 32 - 1 downto 28 * 32) when "11100",
			        bram_do(30 * 32 - 1 downto 29 * 32) when "11101",
			        bram_do(31 * 32 - 1 downto 30 * 32) when "11110",
			        bram_do(32 * 32 - 1 downto 31 * 32) when "11111";
	end block output_controller_31;


	bram_inst : for i in 0 to N_PORTS / 2 - 1 generate

		RAMB16BWER_INST : RAMB16BWER

		generic map (

			-- Configurable data with for ports A and B
			DATA_WIDTH_A => 36,
			DATA_WIDTH_B => 36,

			-- Enable RST capability
			EN_RSTRAM_A => TRUE,
			EN_RSTRAM_B => TRUE,

			-- Reset type
			RSTTYPE => "SYNC",

			-- Optional port output register
			DOA_REG => 0,
			DOB_REG => 0,
			-- Priority given to RAM RST over EN pin (when DO[A|B]_REG = 0)
			RST_PRIORITY_A => "SR",
			RST_PRIORITY_B => "SR",

			-- Initial values on ports
			INIT_A => X"000000000",
			INIT_B => X"000000000",
			INIT_FILE => "NONE",

			-- Warning produced and affected outputs/memory location go unknown
			SIM_COLLISION_CHECK => "ALL",

			-- Simulation device (must be set to "SPARTAN6" for proper simulation behavior
			SIM_DEVICE => "SPARTAN6",

			-- Output value on the DO ports upon the assertion of the syncronous reset signal
			SRVAL_A => X"000000000",
			SRVAL_B => X"000000000",

			-- NO_CHANGE mode: the output latches remain unchanged during a write operation
			WRITE_MODE_A => "READ_FIRST",
			WRITE_MODE_B => "READ_FIRST",

			-- Initial contents of the RAM
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

			-- Parity bits initialization
			INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"

		) port map (

			DOA                  => bram_do((2 * i + 1) * 32 - 1 downto (2 * i + 0) * 32),    -- Output port-A data
			DOB                  => bram_do((2 * i + 2) * 32 - 1 downto (2 * i + 1) * 32),    -- Output port-B data
			DOPA                 => open,                                                     -- We are not using parity bits
			DOPB                 => open,                                                     -- We are not using parity bits
			DIA                  => bram_di((2 * i + 1) * 32 - 1 downto (2 * i + 0) * 32),    -- Input port-A data
			DIB                  => bram_di((2 * i + 2) * 32 - 1 downto (2 * i + 1) * 32),    -- Input port-B data
			DIPA                 => DIP_value,                                                -- Input parity bits always set to 0 (not using them)
			DIPB                 => DIP_value,                                                -- Input parity bits always set to 0 (not using them)
			ADDRA(13 downto 5)   => bram_addr((2 * i + 1) * 9 - 1 downto (2 * i + 0) * 9),    -- Input port-A address
			ADDRA(4 downto 0)    => LOWADDR_value,                                            -- Set low adress bits to 0
			ADDRB(13 downto 5)   => bram_addr((2 * i + 2) * 9 - 1 downto (2 * i + 1) * 9),    -- Input port-B address
			ADDRB(4 downto 0)    => LOWADDR_value,                                            -- Set low adress bits to 0
			CLKA                 => BRAM_CLK,                                                 -- Input port-A clock
			CLKB                 => BRAM_CLK,                                                 -- Input port-B clock
			ENA                  => bram_en(2 * i),                                           -- Input port-A enable
			ENB                  => bram_en(2 * i + 1),                                       -- Input port-B enable
			REGCEA               => REGCE_value,                                              -- Input port-A output register enable
			REGCEB               => REGCE_value,                                              -- Input port-B output register enable
			RSTA                 => RST,                                                      -- Input port-A reset
			RSTB                 => RST,                                                      -- Input port-B reset
			WEA                  => bram_we((2 * i + 1) * 4 - 1 downto (2 * i + 0) * 4),      -- Input port-A write enable
			WEB                  => bram_we((2 * i + 2) * 4 - 1 downto (2 * i + 1) * 4)       -- Input port-B write enable

		);

	end generate bram_inst;


end smem_arch;
